
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);
-- GENERATED BY BC_MEM_PACKER
-- DATE: Fri May 31 13:35:18 2019

	signal mem : ram_t := (

	

		255 =>	x"01010101", -- IMG_16x16_1end_down
		256 =>	x"01020203",
		257 =>	x"04010101",
		258 =>	x"01010101",
		259 =>	x"01010101",
		260 =>	x"01020303",
		261 =>	x"02010101",
		262 =>	x"01010101",
		263 =>	x"01010101",
		264 =>	x"01020302",
		265 =>	x"02010101",
		266 =>	x"01010101",
		267 =>	x"01010101",
		268 =>	x"01020203",
		269 =>	x"02010101",
		270 =>	x"01010101",
		271 =>	x"01010101",
		272 =>	x"01020503",
		273 =>	x"02010101",
		274 =>	x"01010101",
		275 =>	x"01010101",
		276 =>	x"01020203",
		277 =>	x"02010101",
		278 =>	x"01010101",
		279 =>	x"01010101",
		280 =>	x"01020603",
		281 =>	x"02010101",
		282 =>	x"01010101",
		283 =>	x"01010101",
		284 =>	x"01020303",
		285 =>	x"02010101",
		286 =>	x"01010101",
		287 =>	x"01010101",
		288 =>	x"01020303",
		289 =>	x"02010101",
		290 =>	x"01010101",
		291 =>	x"01010101",
		292 =>	x"02020306",
		293 =>	x"02010101",
		294 =>	x"01010101",
		295 =>	x"01010101",
		296 =>	x"02020302",
		297 =>	x"02010101",
		298 =>	x"01010101",
		299 =>	x"01010101",
		300 =>	x"02020303",
		301 =>	x"02010101",
		302 =>	x"01010101",
		303 =>	x"01010101",
		304 =>	x"02020307",
		305 =>	x"02010101",
		306 =>	x"01010101",
		307 =>	x"01010101",
		308 =>	x"08020203",
		309 =>	x"02010101",
		310 =>	x"01010101",
		311 =>	x"01010101",
		312 =>	x"08020303",
		313 =>	x"02010101",
		314 =>	x"01010101",
		315 =>	x"01010101",
		316 =>	x"01020202",
		317 =>	x"02010101",
		318 =>	x"01010101",
		319 =>	x"09000000", -- IMG_16x16_1end_left
		320 =>	x"000A0000",
		321 =>	x"0B0C0000",
		322 =>	x"00000D0E",
		323 =>	x"000A0000",
		324 =>	x"0F101112",
		325 =>	x"13141516",
		326 =>	x"00000000",
		327 =>	x"00000000",
		328 =>	x"00000000",
		329 =>	x"00001718",
		330 =>	x"191A1B1C",
		331 =>	x"00001B1B",
		332 =>	x"1D1E1F20",
		333 =>	x"00000000",
		334 =>	x"00000000",
		335 =>	x"00000000",
		336 =>	x"00000000",
		337 =>	x"00000000",
		338 =>	x"00000000",
		339 =>	x"00000000",
		340 =>	x"00000000",
		341 =>	x"00000000",
		342 =>	x"00000000",
		343 =>	x"00000000",
		344 =>	x"00212223",
		345 =>	x"24252600",
		346 =>	x"00000000",
		347 =>	x"00000000",
		348 =>	x"00000000",
		349 =>	x"00000000",
		350 =>	x"00000000",
		351 =>	x"00000000",
		352 =>	x"00000000",
		353 =>	x"00000000",
		354 =>	x"00000000",
		355 =>	x"00000000",
		356 =>	x"00000000",
		357 =>	x"00000000",
		358 =>	x"00000000",
		359 =>	x"00000000",
		360 =>	x"00000000",
		361 =>	x"00000000",
		362 =>	x"00000000",
		363 =>	x"00000000",
		364 =>	x"00000000",
		365 =>	x"00000000",
		366 =>	x"00000000",
		367 =>	x"27272828",
		368 =>	x"291E2A2B",
		369 =>	x"00000000",
		370 =>	x"00000000",
		371 =>	x"27272727",
		372 =>	x"27272727",
		373 =>	x"27272727",
		374 =>	x"27272727",
		375 =>	x"27272727",
		376 =>	x"27272727",
		377 =>	x"27272727",
		378 =>	x"27272727",
		379 =>	x"2C2D2E2F",
		380 =>	x"301E2A2B",
		381 =>	x"27272727",
		382 =>	x"27272727",
		383 =>	x"09000000", -- IMG_16x16_1end_right
		384 =>	x"000A0000",
		385 =>	x"0B0C0000",
		386 =>	x"00000D0E",
		387 =>	x"000A0000",
		388 =>	x"0F101112",
		389 =>	x"13141516",
		390 =>	x"00000000",
		391 =>	x"00000000",
		392 =>	x"00000000",
		393 =>	x"00001718",
		394 =>	x"191A1B1C",
		395 =>	x"00001B1B",
		396 =>	x"1D1E1F20",
		397 =>	x"00000000",
		398 =>	x"00000000",
		399 =>	x"00000000",
		400 =>	x"00000000",
		401 =>	x"00000000",
		402 =>	x"00000000",
		403 =>	x"00000000",
		404 =>	x"00000000",
		405 =>	x"00000000",
		406 =>	x"00000000",
		407 =>	x"00000000",
		408 =>	x"00212223",
		409 =>	x"24252600",
		410 =>	x"00000000",
		411 =>	x"00000000",
		412 =>	x"00000000",
		413 =>	x"00000000",
		414 =>	x"00000000",
		415 =>	x"00000000",
		416 =>	x"00000000",
		417 =>	x"00000000",
		418 =>	x"00000000",
		419 =>	x"00000000",
		420 =>	x"00000000",
		421 =>	x"00000000",
		422 =>	x"00000000",
		423 =>	x"00000000",
		424 =>	x"00000000",
		425 =>	x"00000000",
		426 =>	x"00000000",
		427 =>	x"00000000",
		428 =>	x"00000000",
		429 =>	x"00000000",
		430 =>	x"00000000",
		431 =>	x"27273128",
		432 =>	x"291E2A2B",
		433 =>	x"00000000",
		434 =>	x"00000000",
		435 =>	x"27272727",
		436 =>	x"27272727",
		437 =>	x"27272727",
		438 =>	x"27272727",
		439 =>	x"27272727",
		440 =>	x"27272727",
		441 =>	x"27272727",
		442 =>	x"27272727",
		443 =>	x"2C2D2E2F",
		444 =>	x"301E2A2B",
		445 =>	x"27272727",
		446 =>	x"27272727",
		447 =>	x"09000000", -- IMG_16x16_1end_up
		448 =>	x"000A0000",
		449 =>	x"0B0C0000",
		450 =>	x"00000D0E",
		451 =>	x"000A0000",
		452 =>	x"0F101112",
		453 =>	x"13141516",
		454 =>	x"00000000",
		455 =>	x"00000000",
		456 =>	x"00000000",
		457 =>	x"00001718",
		458 =>	x"191A1B1C",
		459 =>	x"00001B1B",
		460 =>	x"1D1E1F20",
		461 =>	x"00000000",
		462 =>	x"00000000",
		463 =>	x"00000000",
		464 =>	x"00000000",
		465 =>	x"00000000",
		466 =>	x"00000000",
		467 =>	x"00000000",
		468 =>	x"00000000",
		469 =>	x"00000000",
		470 =>	x"00000000",
		471 =>	x"00000000",
		472 =>	x"00212223",
		473 =>	x"24252600",
		474 =>	x"00000000",
		475 =>	x"00000000",
		476 =>	x"00000000",
		477 =>	x"00000000",
		478 =>	x"00000000",
		479 =>	x"00000000",
		480 =>	x"00000000",
		481 =>	x"00000000",
		482 =>	x"00000000",
		483 =>	x"00000000",
		484 =>	x"00000000",
		485 =>	x"00000000",
		486 =>	x"00000000",
		487 =>	x"00000000",
		488 =>	x"00000000",
		489 =>	x"00000000",
		490 =>	x"00000000",
		491 =>	x"00000000",
		492 =>	x"00000000",
		493 =>	x"00000000",
		494 =>	x"00000000",
		495 =>	x"27273128",
		496 =>	x"291E2A2B",
		497 =>	x"00000000",
		498 =>	x"00000000",
		499 =>	x"27272727",
		500 =>	x"27272727",
		501 =>	x"27272727",
		502 =>	x"27272727",
		503 =>	x"27272727",
		504 =>	x"27272727",
		505 =>	x"27272727",
		506 =>	x"27272727",
		507 =>	x"2C2D2E2F",
		508 =>	x"301E2A2B",
		509 =>	x"27272727",
		510 =>	x"27272727",
		511 =>	x"01010101", -- IMG_16x16_1intersection
		512 =>	x"01010232",
		513 =>	x"06020101",
		514 =>	x"01010101",
		515 =>	x"01010101",
		516 =>	x"01010206",
		517 =>	x"06020101",
		518 =>	x"01010101",
		519 =>	x"01010101",
		520 =>	x"01010206",
		521 =>	x"06020101",
		522 =>	x"01010101",
		523 =>	x"01010101",
		524 =>	x"01020206",
		525 =>	x"06020201",
		526 =>	x"01010101",
		527 =>	x"01010101",
		528 =>	x"02020233",
		529 =>	x"06340201",
		530 =>	x"01010101",
		531 =>	x"01010102",
		532 =>	x"02023533",
		533 =>	x"06333436",
		534 =>	x"36010101",
		535 =>	x"08080204",
		536 =>	x"37380606",
		537 =>	x"06063239",
		538 =>	x"02023A08",
		539 =>	x"3B3B3B3C",
		540 =>	x"06060605",
		541 =>	x"06060606",
		542 =>	x"3D060606",
		543 =>	x"063E0606",
		544 =>	x"06060606",
		545 =>	x"06060606",
		546 =>	x"06060606",
		547 =>	x"3F023F06",
		548 =>	x"40060606",
		549 =>	x"40060640",
		550 =>	x"41020404",
		551 =>	x"01010142",
		552 =>	x"43060633",
		553 =>	x"06064445",
		554 =>	x"46010101",
		555 =>	x"01010101",
		556 =>	x"47480606",
		557 =>	x"3D060449",
		558 =>	x"01010101",
		559 =>	x"01010101",
		560 =>	x"01024A40",
		561 =>	x"404B0201",
		562 =>	x"01010101",
		563 =>	x"01010101",
		564 =>	x"014C024D",
		565 =>	x"4D020101",
		566 =>	x"01010101",
		567 =>	x"01010101",
		568 =>	x"01010206",
		569 =>	x"06020101",
		570 =>	x"01010101",
		571 =>	x"01010101",
		572 =>	x"0101024E",
		573 =>	x"06020101",
		574 =>	x"01010101",
		575 =>	x"01010101", -- IMG_16x16_1middle_horizontal
		576 =>	x"01010101",
		577 =>	x"01010101",
		578 =>	x"01010101",
		579 =>	x"01010101",
		580 =>	x"01010101",
		581 =>	x"01010101",
		582 =>	x"01010101",
		583 =>	x"01010101",
		584 =>	x"01010101",
		585 =>	x"01010101",
		586 =>	x"01010101",
		587 =>	x"01010101",
		588 =>	x"01010101",
		589 =>	x"01010101",
		590 =>	x"01010101",
		591 =>	x"01010101",
		592 =>	x"01010101",
		593 =>	x"01010101",
		594 =>	x"01010101",
		595 =>	x"01010101",
		596 =>	x"01010101",
		597 =>	x"01010101",
		598 =>	x"01010101",
		599 =>	x"024F4F02",
		600 =>	x"02020202",
		601 =>	x"02024F4F",
		602 =>	x"4F4F4F02",
		603 =>	x"50515150",
		604 =>	x"51515151",
		605 =>	x"51515151",
		606 =>	x"51515102",
		607 =>	x"51515151",
		608 =>	x"51515151",
		609 =>	x"51515151",
		610 =>	x"51515151",
		611 =>	x"02515151",
		612 =>	x"51515151",
		613 =>	x"51515151",
		614 =>	x"51515152",
		615 =>	x"02535302",
		616 =>	x"02020202",
		617 =>	x"02020202",
		618 =>	x"02020202",
		619 =>	x"01010101",
		620 =>	x"01010101",
		621 =>	x"01010101",
		622 =>	x"01010101",
		623 =>	x"01010101",
		624 =>	x"01010101",
		625 =>	x"01010101",
		626 =>	x"01010101",
		627 =>	x"01010101",
		628 =>	x"01010101",
		629 =>	x"01010101",
		630 =>	x"01010101",
		631 =>	x"01010101",
		632 =>	x"01010101",
		633 =>	x"01010101",
		634 =>	x"01010101",
		635 =>	x"01010101",
		636 =>	x"01010101",
		637 =>	x"01010101",
		638 =>	x"01010101",
		639 =>	x"09000000", -- IMG_16x16_1middle_vertical
		640 =>	x"000A0000",
		641 =>	x"0B0C0000",
		642 =>	x"00000D0E",
		643 =>	x"000A0000",
		644 =>	x"0F101112",
		645 =>	x"13141516",
		646 =>	x"00000000",
		647 =>	x"00000000",
		648 =>	x"00000000",
		649 =>	x"00001718",
		650 =>	x"191A1B1C",
		651 =>	x"00001B1B",
		652 =>	x"1D1E1F20",
		653 =>	x"00000000",
		654 =>	x"00000000",
		655 =>	x"00000000",
		656 =>	x"00000000",
		657 =>	x"00000000",
		658 =>	x"00000000",
		659 =>	x"00000000",
		660 =>	x"00000000",
		661 =>	x"00000000",
		662 =>	x"00000000",
		663 =>	x"00000000",
		664 =>	x"00212223",
		665 =>	x"24252600",
		666 =>	x"00000000",
		667 =>	x"00000000",
		668 =>	x"00000000",
		669 =>	x"00000000",
		670 =>	x"00000000",
		671 =>	x"00000000",
		672 =>	x"00000000",
		673 =>	x"00000000",
		674 =>	x"00000000",
		675 =>	x"00000000",
		676 =>	x"00000000",
		677 =>	x"00000000",
		678 =>	x"00000000",
		679 =>	x"00000000",
		680 =>	x"00000000",
		681 =>	x"00000000",
		682 =>	x"00000000",
		683 =>	x"00000000",
		684 =>	x"00000000",
		685 =>	x"00000000",
		686 =>	x"00000000",
		687 =>	x"27272727",
		688 =>	x"27272727",
		689 =>	x"54555657",
		690 =>	x"58000000",
		691 =>	x"27272727",
		692 =>	x"27272727",
		693 =>	x"27272727",
		694 =>	x"27272727",
		695 =>	x"27272727",
		696 =>	x"27272727",
		697 =>	x"27272727",
		698 =>	x"27272727",
		699 =>	x"2C2D2E2F",
		700 =>	x"301E2A2B",
		701 =>	x"27272727",
		702 =>	x"27272727",
		703 =>	x"01015902", -- IMG_16x16_2end_down
		704 =>	x"5A5A5A5A",
		705 =>	x"5A355B01",
		706 =>	x"01010101",
		707 =>	x"01015C5B",
		708 =>	x"5A5A5A5A",
		709 =>	x"5A5D5901",
		710 =>	x"01010101",
		711 =>	x"01015C5E",
		712 =>	x"5A5A5A5A",
		713 =>	x"5A5F0101",
		714 =>	x"01010101",
		715 =>	x"01015C02",
		716 =>	x"5A5A5A5A",
		717 =>	x"5A025B01",
		718 =>	x"01010101",
		719 =>	x"01010159",
		720 =>	x"5A5A5A5A",
		721 =>	x"5A605B01",
		722 =>	x"01010101",
		723 =>	x"0101015B",
		724 =>	x"5A5A5A5A",
		725 =>	x"5A355B01",
		726 =>	x"01010101",
		727 =>	x"01015C02",
		728 =>	x"5A5A5A5A",
		729 =>	x"5A025B01",
		730 =>	x"01010101",
		731 =>	x"01015C5E",
		732 =>	x"5A5A5A5A",
		733 =>	x"5A025B01",
		734 =>	x"01010101",
		735 =>	x"01015C5B",
		736 =>	x"5A5A5A5A",
		737 =>	x"5A356101",
		738 =>	x"01010101",
		739 =>	x"01015C5E",
		740 =>	x"5A5A5A5A",
		741 =>	x"5A5D5901",
		742 =>	x"01010101",
		743 =>	x"01015C5B",
		744 =>	x"5A5A5A5A",
		745 =>	x"5A025B01",
		746 =>	x"01010101",
		747 =>	x"0101015B",
		748 =>	x"5A5A5A5A",
		749 =>	x"5A5D5901",
		750 =>	x"01010101",
		751 =>	x"01015C5E",
		752 =>	x"625A5A5A",
		753 =>	x"5A025B01",
		754 =>	x"01010101",
		755 =>	x"0101015B",
		756 =>	x"025A5A5A",
		757 =>	x"635D5901",
		758 =>	x"01010101",
		759 =>	x"0101015B",
		760 =>	x"02020202",
		761 =>	x"5D590101",
		762 =>	x"01010101",
		763 =>	x"01010164",
		764 =>	x"59656667",
		765 =>	x"5B590101",
		766 =>	x"01010101",
		767 =>	x"09000000", -- IMG_16x16_2end_left
		768 =>	x"000A0000",
		769 =>	x"0B0C0000",
		770 =>	x"00000D0E",
		771 =>	x"000A0000",
		772 =>	x"0F101112",
		773 =>	x"13141516",
		774 =>	x"00000000",
		775 =>	x"00000000",
		776 =>	x"00000000",
		777 =>	x"00001718",
		778 =>	x"191A1B1C",
		779 =>	x"00001B1B",
		780 =>	x"1D1E1F20",
		781 =>	x"00000000",
		782 =>	x"00000000",
		783 =>	x"00000000",
		784 =>	x"00000000",
		785 =>	x"00000000",
		786 =>	x"00000000",
		787 =>	x"00000000",
		788 =>	x"00000000",
		789 =>	x"00000000",
		790 =>	x"00000000",
		791 =>	x"00000000",
		792 =>	x"00212223",
		793 =>	x"24252600",
		794 =>	x"00000000",
		795 =>	x"00000000",
		796 =>	x"00000000",
		797 =>	x"00000000",
		798 =>	x"00000000",
		799 =>	x"00000000",
		800 =>	x"00000000",
		801 =>	x"00000000",
		802 =>	x"00000000",
		803 =>	x"00000000",
		804 =>	x"00000000",
		805 =>	x"00000000",
		806 =>	x"00000000",
		807 =>	x"00000000",
		808 =>	x"00000000",
		809 =>	x"00000000",
		810 =>	x"00000000",
		811 =>	x"00000000",
		812 =>	x"00000000",
		813 =>	x"00000000",
		814 =>	x"00000000",
		815 =>	x"27273128",
		816 =>	x"291E2A2B",
		817 =>	x"54555657",
		818 =>	x"58000000",
		819 =>	x"27272727",
		820 =>	x"27272727",
		821 =>	x"27272727",
		822 =>	x"27272727",
		823 =>	x"27272727",
		824 =>	x"27272727",
		825 =>	x"27272727",
		826 =>	x"27272727",
		827 =>	x"2C2D2E2F",
		828 =>	x"301E2A2B",
		829 =>	x"27272727",
		830 =>	x"27272727",
		831 =>	x"09000000", -- IMG_16x16_2end_right
		832 =>	x"000A0000",
		833 =>	x"0B0C0000",
		834 =>	x"00000D0E",
		835 =>	x"000A0000",
		836 =>	x"0F101112",
		837 =>	x"13141516",
		838 =>	x"00000000",
		839 =>	x"00000000",
		840 =>	x"00000000",
		841 =>	x"00001718",
		842 =>	x"191A1B1C",
		843 =>	x"00001B1B",
		844 =>	x"1D1E1F20",
		845 =>	x"00000000",
		846 =>	x"00000000",
		847 =>	x"00000000",
		848 =>	x"00000000",
		849 =>	x"00000000",
		850 =>	x"00000000",
		851 =>	x"00000000",
		852 =>	x"00000000",
		853 =>	x"00000000",
		854 =>	x"00000000",
		855 =>	x"00000000",
		856 =>	x"00212223",
		857 =>	x"24252600",
		858 =>	x"00000000",
		859 =>	x"00000000",
		860 =>	x"00000000",
		861 =>	x"00000000",
		862 =>	x"00000000",
		863 =>	x"00000000",
		864 =>	x"00000000",
		865 =>	x"00000000",
		866 =>	x"00000000",
		867 =>	x"00000000",
		868 =>	x"00000000",
		869 =>	x"00000000",
		870 =>	x"00000000",
		871 =>	x"00000000",
		872 =>	x"00000000",
		873 =>	x"00000000",
		874 =>	x"00000000",
		875 =>	x"00000000",
		876 =>	x"00000000",
		877 =>	x"00000000",
		878 =>	x"00000000",
		879 =>	x"27273128",
		880 =>	x"291E2A2B",
		881 =>	x"54555657",
		882 =>	x"58000000",
		883 =>	x"27272727",
		884 =>	x"27272727",
		885 =>	x"27272727",
		886 =>	x"27272727",
		887 =>	x"27272727",
		888 =>	x"27272727",
		889 =>	x"27272727",
		890 =>	x"27272727",
		891 =>	x"2C2D2E2F",
		892 =>	x"301E2A2B",
		893 =>	x"27272727",
		894 =>	x"27272727",
		895 =>	x"09000000", -- IMG_16x16_2end_up
		896 =>	x"000A0000",
		897 =>	x"0B0C0000",
		898 =>	x"00000D0E",
		899 =>	x"000A0000",
		900 =>	x"0F101112",
		901 =>	x"13141516",
		902 =>	x"00000000",
		903 =>	x"00000000",
		904 =>	x"00000000",
		905 =>	x"00001718",
		906 =>	x"191A1B1C",
		907 =>	x"00001B1B",
		908 =>	x"1D1E1F20",
		909 =>	x"00000000",
		910 =>	x"00000000",
		911 =>	x"00000000",
		912 =>	x"00000000",
		913 =>	x"00000000",
		914 =>	x"00000000",
		915 =>	x"00000000",
		916 =>	x"00000000",
		917 =>	x"00000000",
		918 =>	x"00000000",
		919 =>	x"00000000",
		920 =>	x"00212223",
		921 =>	x"24252600",
		922 =>	x"00000000",
		923 =>	x"00000000",
		924 =>	x"00000000",
		925 =>	x"00000000",
		926 =>	x"00000000",
		927 =>	x"00000000",
		928 =>	x"00000000",
		929 =>	x"00000000",
		930 =>	x"00000000",
		931 =>	x"00000000",
		932 =>	x"00000000",
		933 =>	x"00000000",
		934 =>	x"00000000",
		935 =>	x"00000000",
		936 =>	x"00000000",
		937 =>	x"00000000",
		938 =>	x"00000000",
		939 =>	x"00000000",
		940 =>	x"00000000",
		941 =>	x"00000000",
		942 =>	x"00000000",
		943 =>	x"27273128",
		944 =>	x"291E2A2B",
		945 =>	x"54555657",
		946 =>	x"58000000",
		947 =>	x"27272727",
		948 =>	x"27272727",
		949 =>	x"27272727",
		950 =>	x"27272727",
		951 =>	x"27272727",
		952 =>	x"27272727",
		953 =>	x"27272727",
		954 =>	x"27272727",
		955 =>	x"2C2D2E2F",
		956 =>	x"301E2A2B",
		957 =>	x"27272727",
		958 =>	x"27272727",
		959 =>	x"01010101", -- IMG_16x16_2intersection
		960 =>	x"59026869",
		961 =>	x"696A0259",
		962 =>	x"01010101",
		963 =>	x"01010101",
		964 =>	x"5B026969",
		965 =>	x"69690259",
		966 =>	x"01010101",
		967 =>	x"01010159",
		968 =>	x"02026969",
		969 =>	x"69690259",
		970 =>	x"01010101",
		971 =>	x"0101645E",
		972 =>	x"02696969",
		973 =>	x"69690202",
		974 =>	x"5E640101",
		975 =>	x"6B596502",
		976 =>	x"6C696969",
		977 =>	x"69696902",
		978 =>	x"0265596B",
		979 =>	x"6D026C6C",
		980 =>	x"69696969",
		981 =>	x"6969696E",
		982 =>	x"6F6C026D",
		983 =>	x"70696969",
		984 =>	x"69696969",
		985 =>	x"69696969",
		986 =>	x"69696970",
		987 =>	x"69696969",
		988 =>	x"69696969",
		989 =>	x"69696969",
		990 =>	x"69696969",
		991 =>	x"69696969",
		992 =>	x"69696969",
		993 =>	x"69696969",
		994 =>	x"69696969",
		995 =>	x"69696969",
		996 =>	x"69696969",
		997 =>	x"69696969",
		998 =>	x"69696969",
		999 =>	x"35350269",
		1000 =>	x"69696969",
		1001 =>	x"69696969",
		1002 =>	x"69023535",
		1003 =>	x"715B5D02",
		1004 =>	x"35696969",
		1005 =>	x"69696902",
		1006 =>	x"025D5B71",
		1007 =>	x"0101595D",
		1008 =>	x"02696969",
		1009 =>	x"69696902",
		1010 =>	x"02590101",
		1011 =>	x"01010159",
		1012 =>	x"02696969",
		1013 =>	x"69690272",
		1014 =>	x"5B590101",
		1015 =>	x"01010101",
		1016 =>	x"73696969",
		1017 =>	x"69690259",
		1018 =>	x"59010101",
		1019 =>	x"01010101",
		1020 =>	x"59026A69",
		1021 =>	x"696A7459",
		1022 =>	x"01010101",
		1023 =>	x"01010101", -- IMG_16x16_2middle_horizontal
		1024 =>	x"01010101",
		1025 =>	x"01010101",
		1026 =>	x"01010101",
		1027 =>	x"01010101",
		1028 =>	x"01010101",
		1029 =>	x"01010101",
		1030 =>	x"01010101",
		1031 =>	x"01010101",
		1032 =>	x"01010101",
		1033 =>	x"01010101",
		1034 =>	x"01010101",
		1035 =>	x"01010101",
		1036 =>	x"01010101",
		1037 =>	x"01010101",
		1038 =>	x"01010101",
		1039 =>	x"01010101",
		1040 =>	x"01010101",
		1041 =>	x"01010101",
		1042 =>	x"01010101",
		1043 =>	x"01010101",
		1044 =>	x"01010101",
		1045 =>	x"01010101",
		1046 =>	x"01010101",
		1047 =>	x"02020202",
		1048 =>	x"02020202",
		1049 =>	x"02020202",
		1050 =>	x"02020202",
		1051 =>	x"50510206",
		1052 =>	x"06060606",
		1053 =>	x"06060606",
		1054 =>	x"06060602",
		1055 =>	x"51065106",
		1056 =>	x"06060606",
		1057 =>	x"06065106",
		1058 =>	x"06060606",
		1059 =>	x"02060606",
		1060 =>	x"06060606",
		1061 =>	x"06060606",
		1062 =>	x"06060606",
		1063 =>	x"02020202",
		1064 =>	x"02020202",
		1065 =>	x"02020202",
		1066 =>	x"02020202",
		1067 =>	x"01010101",
		1068 =>	x"01010101",
		1069 =>	x"01010101",
		1070 =>	x"01010101",
		1071 =>	x"01010101",
		1072 =>	x"01010101",
		1073 =>	x"01010101",
		1074 =>	x"01010101",
		1075 =>	x"01010101",
		1076 =>	x"01010101",
		1077 =>	x"01010101",
		1078 =>	x"01010101",
		1079 =>	x"01010101",
		1080 =>	x"01010101",
		1081 =>	x"01010101",
		1082 =>	x"01010101",
		1083 =>	x"01010101",
		1084 =>	x"01010101",
		1085 =>	x"01010101",
		1086 =>	x"01010101",
		1087 =>	x"09000000", -- IMG_16x16_2middle_vertical
		1088 =>	x"000A0000",
		1089 =>	x"0B0C0000",
		1090 =>	x"00000D0E",
		1091 =>	x"000A0000",
		1092 =>	x"0F101112",
		1093 =>	x"13141516",
		1094 =>	x"00000000",
		1095 =>	x"00000000",
		1096 =>	x"00000000",
		1097 =>	x"00001718",
		1098 =>	x"191A1B1C",
		1099 =>	x"00001B1B",
		1100 =>	x"1D1E1F20",
		1101 =>	x"00000000",
		1102 =>	x"00000000",
		1103 =>	x"00000000",
		1104 =>	x"00000000",
		1105 =>	x"00000000",
		1106 =>	x"00000000",
		1107 =>	x"00000000",
		1108 =>	x"00000000",
		1109 =>	x"00000000",
		1110 =>	x"00000000",
		1111 =>	x"00000000",
		1112 =>	x"00212223",
		1113 =>	x"24252600",
		1114 =>	x"00000000",
		1115 =>	x"00000000",
		1116 =>	x"00000000",
		1117 =>	x"00000000",
		1118 =>	x"00000000",
		1119 =>	x"00000000",
		1120 =>	x"00000000",
		1121 =>	x"00000000",
		1122 =>	x"00000000",
		1123 =>	x"00000000",
		1124 =>	x"00000000",
		1125 =>	x"00000000",
		1126 =>	x"00000000",
		1127 =>	x"00000000",
		1128 =>	x"00000000",
		1129 =>	x"00000000",
		1130 =>	x"00000000",
		1131 =>	x"00000000",
		1132 =>	x"00000000",
		1133 =>	x"00000000",
		1134 =>	x"00000000",
		1135 =>	x"27272727",
		1136 =>	x"27272727",
		1137 =>	x"54555657",
		1138 =>	x"58000000",
		1139 =>	x"27272727",
		1140 =>	x"27272727",
		1141 =>	x"27272727",
		1142 =>	x"27272727",
		1143 =>	x"27272727",
		1144 =>	x"27272727",
		1145 =>	x"27272727",
		1146 =>	x"27272727",
		1147 =>	x"2C2D2E2F",
		1148 =>	x"301E2A2B",
		1149 =>	x"27272727",
		1150 =>	x"27272727",
		1151 =>	x"09000000", -- IMG_16x16_3end_down
		1152 =>	x"000A0000",
		1153 =>	x"0B0C0000",
		1154 =>	x"00000D0E",
		1155 =>	x"000A0000",
		1156 =>	x"0F101112",
		1157 =>	x"13141516",
		1158 =>	x"00000000",
		1159 =>	x"00000000",
		1160 =>	x"00000000",
		1161 =>	x"00001718",
		1162 =>	x"191A1B1C",
		1163 =>	x"00001B1B",
		1164 =>	x"1D1E1F20",
		1165 =>	x"00000000",
		1166 =>	x"00000000",
		1167 =>	x"00000000",
		1168 =>	x"00000000",
		1169 =>	x"00000000",
		1170 =>	x"00000000",
		1171 =>	x"00000000",
		1172 =>	x"00000000",
		1173 =>	x"00000000",
		1174 =>	x"00000000",
		1175 =>	x"00000000",
		1176 =>	x"00212223",
		1177 =>	x"24252600",
		1178 =>	x"00000000",
		1179 =>	x"00000000",
		1180 =>	x"00000000",
		1181 =>	x"00000000",
		1182 =>	x"00000000",
		1183 =>	x"00000000",
		1184 =>	x"00000000",
		1185 =>	x"00000000",
		1186 =>	x"00000000",
		1187 =>	x"00000000",
		1188 =>	x"00000000",
		1189 =>	x"00000000",
		1190 =>	x"00000000",
		1191 =>	x"00000000",
		1192 =>	x"00000000",
		1193 =>	x"00000000",
		1194 =>	x"00000000",
		1195 =>	x"00000000",
		1196 =>	x"00000000",
		1197 =>	x"00000000",
		1198 =>	x"00000000",
		1199 =>	x"27273128",
		1200 =>	x"291E2A2B",
		1201 =>	x"54555657",
		1202 =>	x"58000000",
		1203 =>	x"27272727",
		1204 =>	x"27272727",
		1205 =>	x"27272727",
		1206 =>	x"27272727",
		1207 =>	x"27272727",
		1208 =>	x"27272727",
		1209 =>	x"27272727",
		1210 =>	x"27272727",
		1211 =>	x"2C2D2E2F",
		1212 =>	x"301E2A2B",
		1213 =>	x"27272727",
		1214 =>	x"27272727",
		1215 =>	x"09000000", -- IMG_16x16_3end_left
		1216 =>	x"000A0000",
		1217 =>	x"0B0C0000",
		1218 =>	x"00000D0E",
		1219 =>	x"000A0000",
		1220 =>	x"0F101112",
		1221 =>	x"13141516",
		1222 =>	x"00000000",
		1223 =>	x"00000000",
		1224 =>	x"00000000",
		1225 =>	x"00001718",
		1226 =>	x"191A1B1C",
		1227 =>	x"00001B1B",
		1228 =>	x"1D1E1F20",
		1229 =>	x"00000000",
		1230 =>	x"00000000",
		1231 =>	x"00000000",
		1232 =>	x"00000000",
		1233 =>	x"00000000",
		1234 =>	x"00000000",
		1235 =>	x"00000000",
		1236 =>	x"00000000",
		1237 =>	x"00000000",
		1238 =>	x"00000000",
		1239 =>	x"00000000",
		1240 =>	x"00212223",
		1241 =>	x"24252600",
		1242 =>	x"00000000",
		1243 =>	x"00000000",
		1244 =>	x"00000000",
		1245 =>	x"00000000",
		1246 =>	x"00000000",
		1247 =>	x"00000000",
		1248 =>	x"00000000",
		1249 =>	x"00000000",
		1250 =>	x"00000000",
		1251 =>	x"00000000",
		1252 =>	x"00000000",
		1253 =>	x"00000000",
		1254 =>	x"00000000",
		1255 =>	x"00000000",
		1256 =>	x"00000000",
		1257 =>	x"00000000",
		1258 =>	x"00000000",
		1259 =>	x"00000000",
		1260 =>	x"00000000",
		1261 =>	x"00000000",
		1262 =>	x"00000000",
		1263 =>	x"27273128",
		1264 =>	x"291E2A2B",
		1265 =>	x"54555657",
		1266 =>	x"58000000",
		1267 =>	x"27272727",
		1268 =>	x"27272727",
		1269 =>	x"27272727",
		1270 =>	x"27272727",
		1271 =>	x"27272727",
		1272 =>	x"27272727",
		1273 =>	x"27272727",
		1274 =>	x"27272727",
		1275 =>	x"2C2D2E2F",
		1276 =>	x"301E2A2B",
		1277 =>	x"27272727",
		1278 =>	x"27272727",
		1279 =>	x"09000000", -- IMG_16x16_3end_right
		1280 =>	x"000A0000",
		1281 =>	x"0B0C0000",
		1282 =>	x"00000D0E",
		1283 =>	x"000A0000",
		1284 =>	x"0F101112",
		1285 =>	x"13141516",
		1286 =>	x"00000000",
		1287 =>	x"00000000",
		1288 =>	x"00000000",
		1289 =>	x"00001718",
		1290 =>	x"191A1B1C",
		1291 =>	x"00001B1B",
		1292 =>	x"1D1E1F20",
		1293 =>	x"00000000",
		1294 =>	x"00000000",
		1295 =>	x"00000000",
		1296 =>	x"00000000",
		1297 =>	x"00000000",
		1298 =>	x"00000000",
		1299 =>	x"00000000",
		1300 =>	x"00000000",
		1301 =>	x"00000000",
		1302 =>	x"00000000",
		1303 =>	x"00000000",
		1304 =>	x"00212223",
		1305 =>	x"24252600",
		1306 =>	x"00000000",
		1307 =>	x"00000000",
		1308 =>	x"00000000",
		1309 =>	x"00000000",
		1310 =>	x"00000000",
		1311 =>	x"00000000",
		1312 =>	x"00000000",
		1313 =>	x"00000000",
		1314 =>	x"00000000",
		1315 =>	x"00000000",
		1316 =>	x"00000000",
		1317 =>	x"00000000",
		1318 =>	x"00000000",
		1319 =>	x"00000000",
		1320 =>	x"00000000",
		1321 =>	x"00000000",
		1322 =>	x"00000000",
		1323 =>	x"00000000",
		1324 =>	x"00000000",
		1325 =>	x"00000000",
		1326 =>	x"00000000",
		1327 =>	x"27273128",
		1328 =>	x"291E2A2B",
		1329 =>	x"54555657",
		1330 =>	x"58000000",
		1331 =>	x"27272727",
		1332 =>	x"27272727",
		1333 =>	x"27272727",
		1334 =>	x"27272727",
		1335 =>	x"27272727",
		1336 =>	x"27272727",
		1337 =>	x"27272727",
		1338 =>	x"27272727",
		1339 =>	x"2C2D2E2F",
		1340 =>	x"301E2A2B",
		1341 =>	x"27272727",
		1342 =>	x"27272727",
		1343 =>	x"01010101", -- IMG_16x16_3end_up
		1344 =>	x"59595959",
		1345 =>	x"59595959",
		1346 =>	x"59590101",
		1347 =>	x"01010101",
		1348 =>	x"5B02755D",
		1349 =>	x"76590202",
		1350 =>	x"5B597701",
		1351 =>	x"0101015B",
		1352 =>	x"02787878",
		1353 =>	x"78787802",
		1354 =>	x"025B0101",
		1355 =>	x"01010179",
		1356 =>	x"35787878",
		1357 =>	x"78787878",
		1358 =>	x"027A7701",
		1359 =>	x"0101015B",
		1360 =>	x"3578787B",
		1361 =>	x"78787878",
		1362 =>	x"7C5B0101",
		1363 =>	x"01010179",
		1364 =>	x"3578787B",
		1365 =>	x"78787878",
		1366 =>	x"7C5B7701",
		1367 =>	x"0101015B",
		1368 =>	x"0278787D",
		1369 =>	x"78787878",
		1370 =>	x"7E7A7701",
		1371 =>	x"0101015D",
		1372 =>	x"7F787880",
		1373 =>	x"78787878",
		1374 =>	x"7C5B7701",
		1375 =>	x"01010179",
		1376 =>	x"35787878",
		1377 =>	x"78787878",
		1378 =>	x"7C7A7701",
		1379 =>	x"01010179",
		1380 =>	x"02787878",
		1381 =>	x"78787878",
		1382 =>	x"78027701",
		1383 =>	x"01010179",
		1384 =>	x"7F787878",
		1385 =>	x"78787878",
		1386 =>	x"785B0101",
		1387 =>	x"01010179",
		1388 =>	x"81787878",
		1389 =>	x"78787878",
		1390 =>	x"78590101",
		1391 =>	x"01010179",
		1392 =>	x"35787878",
		1393 =>	x"78787878",
		1394 =>	x"02027701",
		1395 =>	x"01010159",
		1396 =>	x"82787878",
		1397 =>	x"78787878",
		1398 =>	x"7C7A7701",
		1399 =>	x"0101015B",
		1400 =>	x"35787878",
		1401 =>	x"78787878",
		1402 =>	x"7C5B7701",
		1403 =>	x"01010179",
		1404 =>	x"7F787878",
		1405 =>	x"78787878",
		1406 =>	x"02025901",
		1407 =>	x"01018359", -- IMG_16x16_3intersection
		1408 =>	x"02696969",
		1409 =>	x"69696906",
		1410 =>	x"76590101",
		1411 =>	x"01015902",
		1412 =>	x"05696969",
		1413 =>	x"69696969",
		1414 =>	x"045B0101",
		1415 =>	x"5C597A02",
		1416 =>	x"69696969",
		1417 =>	x"69696969",
		1418 =>	x"8402595C",
		1419 =>	x"5B7C027C",
		1420 =>	x"69696969",
		1421 =>	x"69696969",
		1422 =>	x"6C02025B",
		1423 =>	x"32328569",
		1424 =>	x"69696969",
		1425 =>	x"69696969",
		1426 =>	x"69696969",
		1427 =>	x"69696969",
		1428 =>	x"69696969",
		1429 =>	x"69696969",
		1430 =>	x"69696969",
		1431 =>	x"69696969",
		1432 =>	x"69696969",
		1433 =>	x"69696969",
		1434 =>	x"69696969",
		1435 =>	x"86876969",
		1436 =>	x"69696969",
		1437 =>	x"69696986",
		1438 =>	x"87698686",
		1439 =>	x"69696969",
		1440 =>	x"69696969",
		1441 =>	x"69696969",
		1442 =>	x"69696969",
		1443 =>	x"69696969",
		1444 =>	x"69696969",
		1445 =>	x"69696969",
		1446 =>	x"69696969",
		1447 =>	x"69696969",
		1448 =>	x"69696969",
		1449 =>	x"69696969",
		1450 =>	x"69696969",
		1451 =>	x"88696969",
		1452 =>	x"69696969",
		1453 =>	x"69696969",
		1454 =>	x"69690688",
		1455 =>	x"5D020235",
		1456 =>	x"8969698A",
		1457 =>	x"69696969",
		1458 =>	x"8B02355D",
		1459 =>	x"59728C02",
		1460 =>	x"02696969",
		1461 =>	x"698A6969",
		1462 =>	x"02027259",
		1463 =>	x"018D5902",
		1464 =>	x"02696969",
		1465 =>	x"69696969",
		1466 =>	x"02738D01",
		1467 =>	x"01015979",
		1468 =>	x"028E6969",
		1469 =>	x"69696969",
		1470 =>	x"8F590101",
		1471 =>	x"01010101", -- IMG_16x16_3middle_horizontal
		1472 =>	x"01010101",
		1473 =>	x"01010101",
		1474 =>	x"01010101",
		1475 =>	x"01010101",
		1476 =>	x"01010101",
		1477 =>	x"01010101",
		1478 =>	x"01010101",
		1479 =>	x"90900101",
		1480 =>	x"01909090",
		1481 =>	x"90019090",
		1482 =>	x"01010190",
		1483 =>	x"91925991",
		1484 =>	x"91919191",
		1485 =>	x"93929192",
		1486 =>	x"91925991",
		1487 =>	x"948F7C80",
		1488 =>	x"80809596",
		1489 =>	x"80808080",
		1490 =>	x"80809794",
		1491 =>	x"80808080",
		1492 =>	x"80808080",
		1493 =>	x"80808080",
		1494 =>	x"80808098",
		1495 =>	x"80808080",
		1496 =>	x"80808080",
		1497 =>	x"80808080",
		1498 =>	x"80808080",
		1499 =>	x"80808080",
		1500 =>	x"80808080",
		1501 =>	x"80808080",
		1502 =>	x"80808080",
		1503 =>	x"80808080",
		1504 =>	x"80808080",
		1505 =>	x"80808080",
		1506 =>	x"80808080",
		1507 =>	x"80808080",
		1508 =>	x"80808080",
		1509 =>	x"80808080",
		1510 =>	x"80808080",
		1511 =>	x"80808080",
		1512 =>	x"80808080",
		1513 =>	x"80808080",
		1514 =>	x"80808080",
		1515 =>	x"80808080",
		1516 =>	x"80808080",
		1517 =>	x"80808080",
		1518 =>	x"80808080",
		1519 =>	x"5D808080",
		1520 =>	x"80808080",
		1521 =>	x"80808080",
		1522 =>	x"80028080",
		1523 =>	x"93929993",
		1524 =>	x"59929399",
		1525 =>	x"92999292",
		1526 =>	x"99929999",
		1527 =>	x"599A9A9A",
		1528 =>	x"01019A9A",
		1529 =>	x"9A9A9A01",
		1530 =>	x"9A010101",
		1531 =>	x"01010101",
		1532 =>	x"01010101",
		1533 =>	x"01010101",
		1534 =>	x"01010101",
		1535 =>	x"09000000", -- IMG_16x16_3middle_vertical
		1536 =>	x"000A0000",
		1537 =>	x"0B0C0000",
		1538 =>	x"00000D0E",
		1539 =>	x"000A0000",
		1540 =>	x"0F101112",
		1541 =>	x"13141516",
		1542 =>	x"00000000",
		1543 =>	x"00000000",
		1544 =>	x"00000000",
		1545 =>	x"00001718",
		1546 =>	x"191A1B1C",
		1547 =>	x"00001B1B",
		1548 =>	x"1D1E1F20",
		1549 =>	x"00000000",
		1550 =>	x"00000000",
		1551 =>	x"00000000",
		1552 =>	x"00000000",
		1553 =>	x"00000000",
		1554 =>	x"00000000",
		1555 =>	x"00000000",
		1556 =>	x"00000000",
		1557 =>	x"00000000",
		1558 =>	x"00000000",
		1559 =>	x"00000000",
		1560 =>	x"00212223",
		1561 =>	x"24252600",
		1562 =>	x"00000000",
		1563 =>	x"00000000",
		1564 =>	x"00000000",
		1565 =>	x"00000000",
		1566 =>	x"00000000",
		1567 =>	x"00000000",
		1568 =>	x"00000000",
		1569 =>	x"00000000",
		1570 =>	x"00000000",
		1571 =>	x"00000000",
		1572 =>	x"00000000",
		1573 =>	x"00000000",
		1574 =>	x"00000000",
		1575 =>	x"00000000",
		1576 =>	x"00000000",
		1577 =>	x"00000000",
		1578 =>	x"00000000",
		1579 =>	x"00000000",
		1580 =>	x"00000000",
		1581 =>	x"00000000",
		1582 =>	x"00000000",
		1583 =>	x"27272727",
		1584 =>	x"27272727",
		1585 =>	x"54555657",
		1586 =>	x"58000000",
		1587 =>	x"27272727",
		1588 =>	x"27272727",
		1589 =>	x"27272727",
		1590 =>	x"27272727",
		1591 =>	x"27272727",
		1592 =>	x"27272727",
		1593 =>	x"27272727",
		1594 =>	x"27272727",
		1595 =>	x"2C2D2E2F",
		1596 =>	x"301E2A2B",
		1597 =>	x"27272727",
		1598 =>	x"27272727",
		1599 =>	x"59027C9B", -- IMG_16x16_4end_down
		1600 =>	x"7B9C9D7B",
		1601 =>	x"7B7B7B9C",
		1602 =>	x"02720101",
		1603 =>	x"835B027B",
		1604 =>	x"7B7B7B7B",
		1605 =>	x"7B7B7B7B",
		1606 =>	x"025B0101",
		1607 =>	x"839E027B",
		1608 =>	x"7B7B7B7B",
		1609 =>	x"7B7B7B7B",
		1610 =>	x"025B0101",
		1611 =>	x"8302027B",
		1612 =>	x"7B7B7B7B",
		1613 =>	x"7B7B7B7B",
		1614 =>	x"02720101",
		1615 =>	x"0159027B",
		1616 =>	x"7B7B7B7B",
		1617 =>	x"7B7B7B7B",
		1618 =>	x"02720101",
		1619 =>	x"015B027B",
		1620 =>	x"7B7B7B7B",
		1621 =>	x"7B7B7B7B",
		1622 =>	x"02720101",
		1623 =>	x"8302027B",
		1624 =>	x"7B7B7B7B",
		1625 =>	x"7B7B7B9F",
		1626 =>	x"02720101",
		1627 =>	x"839E7B7B",
		1628 =>	x"7B7B7B7B",
		1629 =>	x"7B7B7B7B",
		1630 =>	x"02720101",
		1631 =>	x"835BA07B",
		1632 =>	x"7B7B7B7B",
		1633 =>	x"7B7B7B7B",
		1634 =>	x"028C0101",
		1635 =>	x"839E7B7B",
		1636 =>	x"7B7B7B7B",
		1637 =>	x"7B7B7B7B",
		1638 =>	x"02720101",
		1639 =>	x"835BA17B",
		1640 =>	x"7B7B7B7B",
		1641 =>	x"7B7B7B7B",
		1642 =>	x"02720101",
		1643 =>	x"015B7B7B",
		1644 =>	x"7B7B7B7B",
		1645 =>	x"7B7B7B7B",
		1646 =>	x"025B0101",
		1647 =>	x"839E027B",
		1648 =>	x"7B7B7B7B",
		1649 =>	x"7B7B7B35",
		1650 =>	x"02720101",
		1651 =>	x"0159027B",
		1652 =>	x"7B7B7B7B",
		1653 =>	x"7B7B0202",
		1654 =>	x"025B0101",
		1655 =>	x"0177595E",
		1656 =>	x"02020202",
		1657 =>	x"0202025D",
		1658 =>	x"59590101",
		1659 =>	x"01010159",
		1660 =>	x"596D5959",
		1661 =>	x"5959A25B",
		1662 =>	x"01010101",
		1663 =>	x"09000000", -- IMG_16x16_4end_left
		1664 =>	x"000A0000",
		1665 =>	x"0B0C0000",
		1666 =>	x"00000D0E",
		1667 =>	x"000A0000",
		1668 =>	x"0F101112",
		1669 =>	x"13141516",
		1670 =>	x"00000000",
		1671 =>	x"00000000",
		1672 =>	x"00000000",
		1673 =>	x"00001718",
		1674 =>	x"191A1B1C",
		1675 =>	x"00001B1B",
		1676 =>	x"1D1E1F20",
		1677 =>	x"00000000",
		1678 =>	x"00000000",
		1679 =>	x"00000000",
		1680 =>	x"00000000",
		1681 =>	x"00000000",
		1682 =>	x"00000000",
		1683 =>	x"00000000",
		1684 =>	x"00000000",
		1685 =>	x"00000000",
		1686 =>	x"00000000",
		1687 =>	x"00000000",
		1688 =>	x"00212223",
		1689 =>	x"24252600",
		1690 =>	x"00000000",
		1691 =>	x"00000000",
		1692 =>	x"00000000",
		1693 =>	x"00000000",
		1694 =>	x"00000000",
		1695 =>	x"00000000",
		1696 =>	x"00000000",
		1697 =>	x"00000000",
		1698 =>	x"00000000",
		1699 =>	x"00000000",
		1700 =>	x"00000000",
		1701 =>	x"00000000",
		1702 =>	x"00000000",
		1703 =>	x"00000000",
		1704 =>	x"00000000",
		1705 =>	x"00000000",
		1706 =>	x"00000000",
		1707 =>	x"00000000",
		1708 =>	x"00000000",
		1709 =>	x"00000000",
		1710 =>	x"00000000",
		1711 =>	x"27273128",
		1712 =>	x"291E2A2B",
		1713 =>	x"54555657",
		1714 =>	x"58000000",
		1715 =>	x"27272727",
		1716 =>	x"27272727",
		1717 =>	x"27272727",
		1718 =>	x"27272727",
		1719 =>	x"27272727",
		1720 =>	x"27272727",
		1721 =>	x"27272727",
		1722 =>	x"27272727",
		1723 =>	x"2C2D2E2F",
		1724 =>	x"301E2A2B",
		1725 =>	x"27272727",
		1726 =>	x"27272727",
		1727 =>	x"09000000", -- IMG_16x16_4end_right
		1728 =>	x"000A0000",
		1729 =>	x"0B0C0000",
		1730 =>	x"00000D0E",
		1731 =>	x"000A0000",
		1732 =>	x"0F101112",
		1733 =>	x"13141516",
		1734 =>	x"00000000",
		1735 =>	x"00000000",
		1736 =>	x"00000000",
		1737 =>	x"00001718",
		1738 =>	x"191A1B1C",
		1739 =>	x"00001B1B",
		1740 =>	x"1D1E1F20",
		1741 =>	x"00000000",
		1742 =>	x"00000000",
		1743 =>	x"00000000",
		1744 =>	x"00000000",
		1745 =>	x"00000000",
		1746 =>	x"00000000",
		1747 =>	x"00000000",
		1748 =>	x"00000000",
		1749 =>	x"00000000",
		1750 =>	x"00000000",
		1751 =>	x"00000000",
		1752 =>	x"00212223",
		1753 =>	x"24252600",
		1754 =>	x"00000000",
		1755 =>	x"00000000",
		1756 =>	x"00000000",
		1757 =>	x"00000000",
		1758 =>	x"00000000",
		1759 =>	x"00000000",
		1760 =>	x"00000000",
		1761 =>	x"00000000",
		1762 =>	x"00000000",
		1763 =>	x"00000000",
		1764 =>	x"00000000",
		1765 =>	x"00000000",
		1766 =>	x"00000000",
		1767 =>	x"00000000",
		1768 =>	x"00000000",
		1769 =>	x"00000000",
		1770 =>	x"00000000",
		1771 =>	x"00000000",
		1772 =>	x"00000000",
		1773 =>	x"00000000",
		1774 =>	x"00000000",
		1775 =>	x"27273128",
		1776 =>	x"291E2A2B",
		1777 =>	x"54555657",
		1778 =>	x"58000000",
		1779 =>	x"27272727",
		1780 =>	x"27272727",
		1781 =>	x"27272727",
		1782 =>	x"27272727",
		1783 =>	x"27272727",
		1784 =>	x"27272727",
		1785 =>	x"27272727",
		1786 =>	x"27272727",
		1787 =>	x"2C2D2E2F",
		1788 =>	x"301E2A2B",
		1789 =>	x"27272727",
		1790 =>	x"27272727",
		1791 =>	x"09000000", -- IMG_16x16_4end_up
		1792 =>	x"000A0000",
		1793 =>	x"0B0C0000",
		1794 =>	x"00000D0E",
		1795 =>	x"000A0000",
		1796 =>	x"0F101112",
		1797 =>	x"13141516",
		1798 =>	x"00000000",
		1799 =>	x"00000000",
		1800 =>	x"00000000",
		1801 =>	x"00001718",
		1802 =>	x"191A1B1C",
		1803 =>	x"00001B1B",
		1804 =>	x"1D1E1F20",
		1805 =>	x"00000000",
		1806 =>	x"00000000",
		1807 =>	x"00000000",
		1808 =>	x"00000000",
		1809 =>	x"00000000",
		1810 =>	x"00000000",
		1811 =>	x"00000000",
		1812 =>	x"00000000",
		1813 =>	x"00000000",
		1814 =>	x"00000000",
		1815 =>	x"00000000",
		1816 =>	x"00212223",
		1817 =>	x"24252600",
		1818 =>	x"00000000",
		1819 =>	x"00000000",
		1820 =>	x"00000000",
		1821 =>	x"00000000",
		1822 =>	x"00000000",
		1823 =>	x"00000000",
		1824 =>	x"00000000",
		1825 =>	x"00000000",
		1826 =>	x"00000000",
		1827 =>	x"00000000",
		1828 =>	x"00000000",
		1829 =>	x"00000000",
		1830 =>	x"00000000",
		1831 =>	x"00000000",
		1832 =>	x"00000000",
		1833 =>	x"00000000",
		1834 =>	x"00000000",
		1835 =>	x"00000000",
		1836 =>	x"00000000",
		1837 =>	x"00000000",
		1838 =>	x"00000000",
		1839 =>	x"27273128",
		1840 =>	x"291E2A2B",
		1841 =>	x"54555657",
		1842 =>	x"58000000",
		1843 =>	x"27272727",
		1844 =>	x"27272727",
		1845 =>	x"27272727",
		1846 =>	x"27272727",
		1847 =>	x"27272727",
		1848 =>	x"27272727",
		1849 =>	x"27272727",
		1850 =>	x"27272727",
		1851 =>	x"2C2D2E2F",
		1852 =>	x"301E2A2B",
		1853 =>	x"27272727",
		1854 =>	x"27272727",
		1855 =>	x"01835902", -- IMG_16x16_4intersection
		1856 =>	x"A3A49D7B",
		1857 =>	x"7B7B7BA3",
		1858 =>	x"02025901",
		1859 =>	x"77590295",
		1860 =>	x"A57B7B7B",
		1861 =>	x"7B7B7BA5",
		1862 =>	x"A6025977",
		1863 =>	x"5B7A02A7",
		1864 =>	x"7B7B7B7B",
		1865 =>	x"7B7B7B7B",
		1866 =>	x"7BA8A95B",
		1867 =>	x"6C6C6C9C",
		1868 =>	x"7B7B7B7B",
		1869 =>	x"7B7B7B7B",
		1870 =>	x"7B7B9C6C",
		1871 =>	x"A4A57B9D",
		1872 =>	x"7B7B7B7B",
		1873 =>	x"7B7B7B7B",
		1874 =>	x"7B7B7B7B",
		1875 =>	x"9B7B7B7B",
		1876 =>	x"7B7B7B7B",
		1877 =>	x"7B7B7B7B",
		1878 =>	x"7B7B7B7B",
		1879 =>	x"7B7B7B7B",
		1880 =>	x"7B7B7B7B",
		1881 =>	x"7B7B7B7B",
		1882 =>	x"7B7B7B7B",
		1883 =>	x"7B7B7B7B",
		1884 =>	x"7B7B7B7B",
		1885 =>	x"7B7B7B7B",
		1886 =>	x"7B7B7B7B",
		1887 =>	x"7B7B7B7B",
		1888 =>	x"7B7B7B7B",
		1889 =>	x"7B7B7B7B",
		1890 =>	x"7B7B7B7B",
		1891 =>	x"7B7B7B7B",
		1892 =>	x"7B7B7B7B",
		1893 =>	x"7B7B7B7B",
		1894 =>	x"7B7B7B7B",
		1895 =>	x"7B7B7B7B",
		1896 =>	x"7B7B7B7B",
		1897 =>	x"7B7B7B7B",
		1898 =>	x"7B7B7B7B",
		1899 =>	x"AA7B7B7B",
		1900 =>	x"7B7B7B7B",
		1901 =>	x"7B7B7B7B",
		1902 =>	x"7B7B7B7B",
		1903 =>	x"ABAC7B7B",
		1904 =>	x"7B7B7B7B",
		1905 =>	x"7B7B7B7B",
		1906 =>	x"7B7BADAB",
		1907 =>	x"8C8CAE7B",
		1908 =>	x"7B7B7B7B",
		1909 =>	x"7B7B7B7B",
		1910 =>	x"7BAF8C8C",
		1911 =>	x"5959026C",
		1912 =>	x"B07B7B7B",
		1913 =>	x"7B7B7B7B",
		1914 =>	x"7B025959",
		1915 =>	x"0159B102",
		1916 =>	x"9B7B7B7B",
		1917 =>	x"7B7B7B7B",
		1918 =>	x"7B025901",
		1919 =>	x"01010101", -- IMG_16x16_4middle_horizontal
		1920 =>	x"01010101",
		1921 =>	x"01010101",
		1922 =>	x"01010101",
		1923 =>	x"9A9A0101",
		1924 =>	x"019A9A9A",
		1925 =>	x"9A019A9A",
		1926 =>	x"0101019A",
		1927 =>	x"99929299",
		1928 =>	x"99999999",
		1929 =>	x"93999992",
		1930 =>	x"99929299",
		1931 =>	x"02020202",
		1932 =>	x"02020202",
		1933 =>	x"02020202",
		1934 =>	x"028F0202",
		1935 =>	x"B27EA3A3",
		1936 =>	x"7EA3A3A3",
		1937 =>	x"A3A3A3B3",
		1938 =>	x"B4A3B4B4",
		1939 =>	x"A3A3A3A3",
		1940 =>	x"A3A3A3A3",
		1941 =>	x"A3A3A3A3",
		1942 =>	x"A3A3A3A3",
		1943 =>	x"A3A3A3A3",
		1944 =>	x"A3A3A3A3",
		1945 =>	x"A3A3A3A3",
		1946 =>	x"A3A3A3A3",
		1947 =>	x"A3A3A3A3",
		1948 =>	x"A3A3A3A3",
		1949 =>	x"A3A3A3A3",
		1950 =>	x"A3A3A3A3",
		1951 =>	x"A3A3A3A3",
		1952 =>	x"A3A3A3A3",
		1953 =>	x"A3A3A3A3",
		1954 =>	x"A3A3A3A3",
		1955 =>	x"B5A3A3A3",
		1956 =>	x"A3A3A3A3",
		1957 =>	x"A3A3A3A3",
		1958 =>	x"A3A3A3A3",
		1959 =>	x"A3A3A3A3",
		1960 =>	x"A3A3A3A3",
		1961 =>	x"A3A3A3A3",
		1962 =>	x"A3A3A3A3",
		1963 =>	x"A3A3A3A3",
		1964 =>	x"A3A3A3A3",
		1965 =>	x"A3A3A3A3",
		1966 =>	x"A3A3B6A3",
		1967 =>	x"A3A3A3A3",
		1968 =>	x"A3A3A3A3",
		1969 =>	x"A3A3A3A3",
		1970 =>	x"A3A302B7",
		1971 =>	x"B8A3A3A3",
		1972 =>	x"A3A3B902",
		1973 =>	x"BAA3A3A3",
		1974 =>	x"A3B90202",
		1975 =>	x"8292BB82",
		1976 =>	x"599282BB",
		1977 =>	x"92BB9292",
		1978 =>	x"BB92BBBB",
		1979 =>	x"59BCBCBC",
		1980 =>	x"0101BCBC",
		1981 =>	x"BCBCBC01",
		1982 =>	x"BC010101",
		1983 =>	x"09000000", -- IMG_16x16_4middle_vertical
		1984 =>	x"000A0000",
		1985 =>	x"0B0C0000",
		1986 =>	x"00000D0E",
		1987 =>	x"000A0000",
		1988 =>	x"0F101112",
		1989 =>	x"13141516",
		1990 =>	x"00000000",
		1991 =>	x"00000000",
		1992 =>	x"00000000",
		1993 =>	x"00001718",
		1994 =>	x"191A1B1C",
		1995 =>	x"00001B1B",
		1996 =>	x"1D1E1F20",
		1997 =>	x"00000000",
		1998 =>	x"00000000",
		1999 =>	x"00000000",
		2000 =>	x"00000000",
		2001 =>	x"00000000",
		2002 =>	x"00000000",
		2003 =>	x"00000000",
		2004 =>	x"00000000",
		2005 =>	x"00000000",
		2006 =>	x"00000000",
		2007 =>	x"00000000",
		2008 =>	x"00212223",
		2009 =>	x"24252600",
		2010 =>	x"00000000",
		2011 =>	x"00000000",
		2012 =>	x"00000000",
		2013 =>	x"00000000",
		2014 =>	x"00000000",
		2015 =>	x"00000000",
		2016 =>	x"00000000",
		2017 =>	x"00000000",
		2018 =>	x"00000000",
		2019 =>	x"00000000",
		2020 =>	x"00000000",
		2021 =>	x"00000000",
		2022 =>	x"00000000",
		2023 =>	x"00000000",
		2024 =>	x"00000000",
		2025 =>	x"00000000",
		2026 =>	x"00000000",
		2027 =>	x"00000000",
		2028 =>	x"00000000",
		2029 =>	x"00000000",
		2030 =>	x"00000000",
		2031 =>	x"27272727",
		2032 =>	x"27272727",
		2033 =>	x"54555657",
		2034 =>	x"58000000",
		2035 =>	x"27272727",
		2036 =>	x"27272727",
		2037 =>	x"27272727",
		2038 =>	x"27272727",
		2039 =>	x"27272727",
		2040 =>	x"27272727",
		2041 =>	x"27272727",
		2042 =>	x"27272727",
		2043 =>	x"2C2D2E2F",
		2044 =>	x"301E2A2B",
		2045 =>	x"27272727",
		2046 =>	x"27272727",
		2047 =>	x"83595B02", -- IMG_16x16_5end_down
		2048 =>	x"0632BD06",
		2049 =>	x"BE063302",
		2050 =>	x"79590101",
		2051 =>	x"01595B7C",
		2052 =>	x"06BF0606",
		2053 =>	x"06060602",
		2054 =>	x"79590101",
		2055 =>	x"0159597C",
		2056 =>	x"06060606",
		2057 =>	x"0606065D",
		2058 =>	x"59C00101",
		2059 =>	x"01595902",
		2060 =>	x"06060606",
		2061 =>	x"0606065D",
		2062 =>	x"59590101",
		2063 =>	x"0159595E",
		2064 =>	x"06060606",
		2065 =>	x"0606BEC1",
		2066 =>	x"79590101",
		2067 =>	x"01595902",
		2068 =>	x"06060606",
		2069 =>	x"06060633",
		2070 =>	x"79590101",
		2071 =>	x"83595902",
		2072 =>	x"06060606",
		2073 =>	x"06060606",
		2074 =>	x"59590101",
		2075 =>	x"0159595E",
		2076 =>	x"06060606",
		2077 =>	x"060606C2",
		2078 =>	x"59590101",
		2079 =>	x"01595902",
		2080 =>	x"06060606",
		2081 =>	x"06060602",
		2082 =>	x"5B590101",
		2083 =>	x"01597A02",
		2084 =>	x"06060606",
		2085 =>	x"06060671",
		2086 =>	x"59590101",
		2087 =>	x"01597A02",
		2088 =>	x"06060606",
		2089 =>	x"0606065B",
		2090 =>	x"59590101",
		2091 =>	x"0159595E",
		2092 =>	x"3D060606",
		2093 =>	x"06060602",
		2094 =>	x"5B590101",
		2095 =>	x"01595B02",
		2096 =>	x"43060606",
		2097 =>	x"0606065D",
		2098 =>	x"59590101",
		2099 =>	x"01595902",
		2100 =>	x"02020202",
		2101 =>	x"4306945B",
		2102 =>	x"59590101",
		2103 =>	x"0101595B",
		2104 =>	x"02020202",
		2105 =>	x"02025D59",
		2106 =>	x"59010101",
		2107 =>	x"0101C364",
		2108 =>	x"C4595959",
		2109 =>	x"765B59C5",
		2110 =>	x"01010101",
		2111 =>	x"09000000", -- IMG_16x16_5end_left
		2112 =>	x"000A0000",
		2113 =>	x"0B0C0000",
		2114 =>	x"00000D0E",
		2115 =>	x"000A0000",
		2116 =>	x"0F101112",
		2117 =>	x"13141516",
		2118 =>	x"00000000",
		2119 =>	x"00000000",
		2120 =>	x"00000000",
		2121 =>	x"00001718",
		2122 =>	x"191A1B1C",
		2123 =>	x"00001B1B",
		2124 =>	x"1D1E1F20",
		2125 =>	x"00000000",
		2126 =>	x"00000000",
		2127 =>	x"00000000",
		2128 =>	x"00000000",
		2129 =>	x"00000000",
		2130 =>	x"00000000",
		2131 =>	x"00000000",
		2132 =>	x"00000000",
		2133 =>	x"00000000",
		2134 =>	x"00000000",
		2135 =>	x"00000000",
		2136 =>	x"00212223",
		2137 =>	x"24252600",
		2138 =>	x"00000000",
		2139 =>	x"00000000",
		2140 =>	x"00000000",
		2141 =>	x"00000000",
		2142 =>	x"00000000",
		2143 =>	x"00000000",
		2144 =>	x"00000000",
		2145 =>	x"00000000",
		2146 =>	x"00000000",
		2147 =>	x"00000000",
		2148 =>	x"00000000",
		2149 =>	x"00000000",
		2150 =>	x"00000000",
		2151 =>	x"00000000",
		2152 =>	x"00000000",
		2153 =>	x"00000000",
		2154 =>	x"00000000",
		2155 =>	x"00000000",
		2156 =>	x"00000000",
		2157 =>	x"00000000",
		2158 =>	x"00000000",
		2159 =>	x"27273128",
		2160 =>	x"291E2A2B",
		2161 =>	x"54555657",
		2162 =>	x"58000000",
		2163 =>	x"27272727",
		2164 =>	x"27272727",
		2165 =>	x"27272727",
		2166 =>	x"27272727",
		2167 =>	x"27272727",
		2168 =>	x"27272727",
		2169 =>	x"27272727",
		2170 =>	x"27272727",
		2171 =>	x"2C2D2E2F",
		2172 =>	x"301E2A2B",
		2173 =>	x"27272727",
		2174 =>	x"27272727",
		2175 =>	x"09000000", -- IMG_16x16_5end_right
		2176 =>	x"000A0000",
		2177 =>	x"0B0C0000",
		2178 =>	x"00000D0E",
		2179 =>	x"000A0000",
		2180 =>	x"0F101112",
		2181 =>	x"13141516",
		2182 =>	x"00000000",
		2183 =>	x"00000000",
		2184 =>	x"00000000",
		2185 =>	x"00001718",
		2186 =>	x"191A1B1C",
		2187 =>	x"00001B1B",
		2188 =>	x"1D1E1F20",
		2189 =>	x"00000000",
		2190 =>	x"00000000",
		2191 =>	x"00000000",
		2192 =>	x"00000000",
		2193 =>	x"00000000",
		2194 =>	x"00000000",
		2195 =>	x"00000000",
		2196 =>	x"00000000",
		2197 =>	x"00000000",
		2198 =>	x"00000000",
		2199 =>	x"00000000",
		2200 =>	x"00212223",
		2201 =>	x"24252600",
		2202 =>	x"00000000",
		2203 =>	x"00000000",
		2204 =>	x"00000000",
		2205 =>	x"00000000",
		2206 =>	x"00000000",
		2207 =>	x"00000000",
		2208 =>	x"00000000",
		2209 =>	x"00000000",
		2210 =>	x"00000000",
		2211 =>	x"00000000",
		2212 =>	x"00000000",
		2213 =>	x"00000000",
		2214 =>	x"00000000",
		2215 =>	x"00000000",
		2216 =>	x"00000000",
		2217 =>	x"00000000",
		2218 =>	x"00000000",
		2219 =>	x"00000000",
		2220 =>	x"00000000",
		2221 =>	x"00000000",
		2222 =>	x"00000000",
		2223 =>	x"27273128",
		2224 =>	x"291E2A2B",
		2225 =>	x"54555657",
		2226 =>	x"58000000",
		2227 =>	x"27272727",
		2228 =>	x"27272727",
		2229 =>	x"27272727",
		2230 =>	x"27272727",
		2231 =>	x"27272727",
		2232 =>	x"27272727",
		2233 =>	x"27272727",
		2234 =>	x"27272727",
		2235 =>	x"2C2D2E2F",
		2236 =>	x"301E2A2B",
		2237 =>	x"27272727",
		2238 =>	x"27272727",
		2239 =>	x"09000000", -- IMG_16x16_5end_up
		2240 =>	x"000A0000",
		2241 =>	x"0B0C0000",
		2242 =>	x"00000D0E",
		2243 =>	x"000A0000",
		2244 =>	x"0F101112",
		2245 =>	x"13141516",
		2246 =>	x"00000000",
		2247 =>	x"00000000",
		2248 =>	x"00000000",
		2249 =>	x"00001718",
		2250 =>	x"191A1B1C",
		2251 =>	x"00001B1B",
		2252 =>	x"1D1E1F20",
		2253 =>	x"00000000",
		2254 =>	x"00000000",
		2255 =>	x"00000000",
		2256 =>	x"00000000",
		2257 =>	x"00000000",
		2258 =>	x"00000000",
		2259 =>	x"00000000",
		2260 =>	x"00000000",
		2261 =>	x"00000000",
		2262 =>	x"00000000",
		2263 =>	x"00000000",
		2264 =>	x"00212223",
		2265 =>	x"24252600",
		2266 =>	x"00000000",
		2267 =>	x"00000000",
		2268 =>	x"00000000",
		2269 =>	x"00000000",
		2270 =>	x"00000000",
		2271 =>	x"00000000",
		2272 =>	x"00000000",
		2273 =>	x"00000000",
		2274 =>	x"00000000",
		2275 =>	x"00000000",
		2276 =>	x"00000000",
		2277 =>	x"00000000",
		2278 =>	x"00000000",
		2279 =>	x"00000000",
		2280 =>	x"00000000",
		2281 =>	x"00000000",
		2282 =>	x"00000000",
		2283 =>	x"00000000",
		2284 =>	x"00000000",
		2285 =>	x"00000000",
		2286 =>	x"00000000",
		2287 =>	x"27273128",
		2288 =>	x"291E2A2B",
		2289 =>	x"54555657",
		2290 =>	x"58000000",
		2291 =>	x"27272727",
		2292 =>	x"27272727",
		2293 =>	x"27272727",
		2294 =>	x"27272727",
		2295 =>	x"27272727",
		2296 =>	x"27272727",
		2297 =>	x"27272727",
		2298 =>	x"27272727",
		2299 =>	x"2C2D2E2F",
		2300 =>	x"301E2A2B",
		2301 =>	x"27272727",
		2302 =>	x"27272727",
		2303 =>	x"01835902", -- IMG_16x16_5intersection
		2304 =>	x"06060606",
		2305 =>	x"06060602",
		2306 =>	x"02590101",
		2307 =>	x"01595902",
		2308 =>	x"C6060606",
		2309 =>	x"06060606",
		2310 =>	x"02595901",
		2311 =>	x"59595902",
		2312 =>	x"06060606",
		2313 =>	x"06060606",
		2314 =>	x"025B5959",
		2315 =>	x"5E020202",
		2316 =>	x"06060606",
		2317 =>	x"06060606",
		2318 =>	x"0202025E",
		2319 =>	x"02020202",
		2320 =>	x"06060606",
		2321 =>	x"06060606",
		2322 =>	x"02020202",
		2323 =>	x"BE6F6F6F",
		2324 =>	x"06060606",
		2325 =>	x"06060606",
		2326 =>	x"BE6F6FBE",
		2327 =>	x"C70606C7",
		2328 =>	x"C7BF0606",
		2329 =>	x"06060606",
		2330 =>	x"06060606",
		2331 =>	x"BD060606",
		2332 =>	x"06060606",
		2333 =>	x"06060606",
		2334 =>	x"06060606",
		2335 =>	x"06060606",
		2336 =>	x"06060606",
		2337 =>	x"06060606",
		2338 =>	x"06060606",
		2339 =>	x"06060606",
		2340 =>	x"06060606",
		2341 =>	x"06060606",
		2342 =>	x"06060606",
		2343 =>	x"C8060606",
		2344 =>	x"06060606",
		2345 =>	x"060606C9",
		2346 =>	x"06060606",
		2347 =>	x"817F8106",
		2348 =>	x"060606BE",
		2349 =>	x"06060606",
		2350 =>	x"CA0606CB",
		2351 =>	x"5D0202BE",
		2352 =>	x"06060606",
		2353 =>	x"06060606",
		2354 =>	x"025D5D5D",
		2355 =>	x"595B0233",
		2356 =>	x"06060606",
		2357 =>	x"06060606",
		2358 =>	x"02595959",
		2359 =>	x"59595B06",
		2360 =>	x"06060606",
		2361 =>	x"06060602",
		2362 =>	x"02595959",
		2363 =>	x"01595902",
		2364 =>	x"06060606",
		2365 =>	x"06060602",
		2366 =>	x"8C590101",
		2367 =>	x"01010101", -- IMG_16x16_5middle_horizontal
		2368 =>	x"01010101",
		2369 =>	x"01010101",
		2370 =>	x"01010101",
		2371 =>	x"01010101",
		2372 =>	x"01010101",
		2373 =>	x"01010101",
		2374 =>	x"01010101",
		2375 =>	x"59599059",
		2376 =>	x"59595959",
		2377 =>	x"59595959",
		2378 =>	x"59599059",
		2379 =>	x"91CC0606",
		2380 =>	x"CD065959",
		2381 =>	x"92595992",
		2382 =>	x"59595992",
		2383 =>	x"CE620606",
		2384 =>	x"0606CF93",
		2385 =>	x"02CF9202",
		2386 =>	x"93929202",
		2387 =>	x"D0060606",
		2388 =>	x"06060606",
		2389 =>	x"06060606",
		2390 =>	x"06060606",
		2391 =>	x"06060606",
		2392 =>	x"06060606",
		2393 =>	x"06060606",
		2394 =>	x"06060606",
		2395 =>	x"06060606",
		2396 =>	x"06060606",
		2397 =>	x"06060606",
		2398 =>	x"06060606",
		2399 =>	x"06060606",
		2400 =>	x"06060606",
		2401 =>	x"06060606",
		2402 =>	x"06060606",
		2403 =>	x"06060606",
		2404 =>	x"06060606",
		2405 =>	x"06060606",
		2406 =>	x"06060606",
		2407 =>	x"06060606",
		2408 =>	x"06060606",
		2409 =>	x"06060606",
		2410 =>	x"06060606",
		2411 =>	x"BE060606",
		2412 =>	x"06060606",
		2413 =>	x"06060606",
		2414 =>	x"06060606",
		2415 =>	x"43060606",
		2416 =>	x"06060606",
		2417 =>	x"06060606",
		2418 =>	x"06060606",
		2419 =>	x"92925959",
		2420 =>	x"59595959",
		2421 =>	x"59999959",
		2422 =>	x"92595959",
		2423 =>	x"59595959",
		2424 =>	x"59595959",
		2425 =>	x"59595959",
		2426 =>	x"59595959",
		2427 =>	x"BC010101",
		2428 =>	x"0101BC01",
		2429 =>	x"01010101",
		2430 =>	x"01010101",
		2431 =>	x"09000000", -- IMG_16x16_5middle_vertical
		2432 =>	x"000A0000",
		2433 =>	x"0B0C0000",
		2434 =>	x"00000D0E",
		2435 =>	x"000A0000",
		2436 =>	x"0F101112",
		2437 =>	x"13141516",
		2438 =>	x"00000000",
		2439 =>	x"00000000",
		2440 =>	x"00000000",
		2441 =>	x"00001718",
		2442 =>	x"191A1B1C",
		2443 =>	x"00001B1B",
		2444 =>	x"1D1E1F20",
		2445 =>	x"00000000",
		2446 =>	x"00000000",
		2447 =>	x"00000000",
		2448 =>	x"00000000",
		2449 =>	x"00000000",
		2450 =>	x"00000000",
		2451 =>	x"00000000",
		2452 =>	x"00000000",
		2453 =>	x"00000000",
		2454 =>	x"00000000",
		2455 =>	x"00000000",
		2456 =>	x"00212223",
		2457 =>	x"24252600",
		2458 =>	x"00000000",
		2459 =>	x"00000000",
		2460 =>	x"00000000",
		2461 =>	x"00000000",
		2462 =>	x"00000000",
		2463 =>	x"00000000",
		2464 =>	x"00000000",
		2465 =>	x"00000000",
		2466 =>	x"00000000",
		2467 =>	x"00000000",
		2468 =>	x"00000000",
		2469 =>	x"00000000",
		2470 =>	x"00000000",
		2471 =>	x"00000000",
		2472 =>	x"00000000",
		2473 =>	x"00000000",
		2474 =>	x"00000000",
		2475 =>	x"00000000",
		2476 =>	x"00000000",
		2477 =>	x"00000000",
		2478 =>	x"00000000",
		2479 =>	x"27272727",
		2480 =>	x"27272727",
		2481 =>	x"54555657",
		2482 =>	x"58000000",
		2483 =>	x"27272727",
		2484 =>	x"27272727",
		2485 =>	x"27272727",
		2486 =>	x"27272727",
		2487 =>	x"27272727",
		2488 =>	x"27272727",
		2489 =>	x"27272727",
		2490 =>	x"27272727",
		2491 =>	x"2C2D2E2F",
		2492 =>	x"301E2A2B",
		2493 =>	x"27272727",
		2494 =>	x"27272727",
		2495 =>	x"09000000", -- IMG_16x16_6end_down
		2496 =>	x"000A0000",
		2497 =>	x"0B0C0000",
		2498 =>	x"00000D0E",
		2499 =>	x"000A0000",
		2500 =>	x"0F101112",
		2501 =>	x"13141516",
		2502 =>	x"00000000",
		2503 =>	x"00000000",
		2504 =>	x"00000000",
		2505 =>	x"00001718",
		2506 =>	x"191A1B1C",
		2507 =>	x"00001B1B",
		2508 =>	x"1D1E1F20",
		2509 =>	x"00000000",
		2510 =>	x"00000000",
		2511 =>	x"00000000",
		2512 =>	x"00000000",
		2513 =>	x"00000000",
		2514 =>	x"00000000",
		2515 =>	x"00000000",
		2516 =>	x"00000000",
		2517 =>	x"00000000",
		2518 =>	x"00000000",
		2519 =>	x"00000000",
		2520 =>	x"00212223",
		2521 =>	x"24252600",
		2522 =>	x"00000000",
		2523 =>	x"00000000",
		2524 =>	x"00000000",
		2525 =>	x"00000000",
		2526 =>	x"00000000",
		2527 =>	x"00000000",
		2528 =>	x"00000000",
		2529 =>	x"00000000",
		2530 =>	x"00000000",
		2531 =>	x"00000000",
		2532 =>	x"00000000",
		2533 =>	x"00000000",
		2534 =>	x"00000000",
		2535 =>	x"00000000",
		2536 =>	x"00000000",
		2537 =>	x"00000000",
		2538 =>	x"00000000",
		2539 =>	x"00000000",
		2540 =>	x"00000000",
		2541 =>	x"00000000",
		2542 =>	x"00000000",
		2543 =>	x"27273128",
		2544 =>	x"291E2A2B",
		2545 =>	x"54555657",
		2546 =>	x"58000000",
		2547 =>	x"27272727",
		2548 =>	x"27272727",
		2549 =>	x"27272727",
		2550 =>	x"27272727",
		2551 =>	x"27272727",
		2552 =>	x"27272727",
		2553 =>	x"27272727",
		2554 =>	x"27272727",
		2555 =>	x"2C2D2E2F",
		2556 =>	x"301E2A2B",
		2557 =>	x"27272727",
		2558 =>	x"27272727",
		2559 =>	x"09000000", -- IMG_16x16_6end_left
		2560 =>	x"000A0000",
		2561 =>	x"0B0C0000",
		2562 =>	x"00000D0E",
		2563 =>	x"000A0000",
		2564 =>	x"0F101112",
		2565 =>	x"13141516",
		2566 =>	x"00000000",
		2567 =>	x"00000000",
		2568 =>	x"00000000",
		2569 =>	x"00001718",
		2570 =>	x"191A1B1C",
		2571 =>	x"00001B1B",
		2572 =>	x"1D1E1F20",
		2573 =>	x"00000000",
		2574 =>	x"00000000",
		2575 =>	x"00000000",
		2576 =>	x"00000000",
		2577 =>	x"00000000",
		2578 =>	x"00000000",
		2579 =>	x"00000000",
		2580 =>	x"00000000",
		2581 =>	x"00000000",
		2582 =>	x"00000000",
		2583 =>	x"00000000",
		2584 =>	x"00212223",
		2585 =>	x"24252600",
		2586 =>	x"00000000",
		2587 =>	x"00000000",
		2588 =>	x"00000000",
		2589 =>	x"00000000",
		2590 =>	x"00000000",
		2591 =>	x"00000000",
		2592 =>	x"00000000",
		2593 =>	x"00000000",
		2594 =>	x"00000000",
		2595 =>	x"00000000",
		2596 =>	x"00000000",
		2597 =>	x"00000000",
		2598 =>	x"00000000",
		2599 =>	x"00000000",
		2600 =>	x"00000000",
		2601 =>	x"00000000",
		2602 =>	x"00000000",
		2603 =>	x"00000000",
		2604 =>	x"00000000",
		2605 =>	x"00000000",
		2606 =>	x"00000000",
		2607 =>	x"27273128",
		2608 =>	x"291E2A2B",
		2609 =>	x"54555657",
		2610 =>	x"58000000",
		2611 =>	x"27272727",
		2612 =>	x"27272727",
		2613 =>	x"27272727",
		2614 =>	x"27272727",
		2615 =>	x"27272727",
		2616 =>	x"27272727",
		2617 =>	x"27272727",
		2618 =>	x"27272727",
		2619 =>	x"2C2D2E2F",
		2620 =>	x"301E2A2B",
		2621 =>	x"27272727",
		2622 =>	x"27272727",
		2623 =>	x"09000000", -- IMG_16x16_6end_right
		2624 =>	x"000A0000",
		2625 =>	x"0B0C0000",
		2626 =>	x"00000D0E",
		2627 =>	x"000A0000",
		2628 =>	x"0F101112",
		2629 =>	x"13141516",
		2630 =>	x"00000000",
		2631 =>	x"00000000",
		2632 =>	x"00000000",
		2633 =>	x"00001718",
		2634 =>	x"191A1B1C",
		2635 =>	x"00001B1B",
		2636 =>	x"1D1E1F20",
		2637 =>	x"00000000",
		2638 =>	x"00000000",
		2639 =>	x"00000000",
		2640 =>	x"00000000",
		2641 =>	x"00000000",
		2642 =>	x"00000000",
		2643 =>	x"00000000",
		2644 =>	x"00000000",
		2645 =>	x"00000000",
		2646 =>	x"00000000",
		2647 =>	x"00000000",
		2648 =>	x"00212223",
		2649 =>	x"24252600",
		2650 =>	x"00000000",
		2651 =>	x"00000000",
		2652 =>	x"00000000",
		2653 =>	x"00000000",
		2654 =>	x"00000000",
		2655 =>	x"00000000",
		2656 =>	x"00000000",
		2657 =>	x"00000000",
		2658 =>	x"00000000",
		2659 =>	x"00000000",
		2660 =>	x"00000000",
		2661 =>	x"00000000",
		2662 =>	x"00000000",
		2663 =>	x"00000000",
		2664 =>	x"00000000",
		2665 =>	x"00000000",
		2666 =>	x"00000000",
		2667 =>	x"00000000",
		2668 =>	x"00000000",
		2669 =>	x"00000000",
		2670 =>	x"00000000",
		2671 =>	x"27273128",
		2672 =>	x"291E2A2B",
		2673 =>	x"54555657",
		2674 =>	x"58000000",
		2675 =>	x"27272727",
		2676 =>	x"27272727",
		2677 =>	x"27272727",
		2678 =>	x"27272727",
		2679 =>	x"27272727",
		2680 =>	x"27272727",
		2681 =>	x"27272727",
		2682 =>	x"27272727",
		2683 =>	x"2C2D2E2F",
		2684 =>	x"301E2A2B",
		2685 =>	x"27272727",
		2686 =>	x"27272727",
		2687 =>	x"01015C59", -- IMG_16x16_6end_up
		2688 =>	x"65D1D2D2",
		2689 =>	x"D2D35D59",
		2690 =>	x"D4010101",
		2691 =>	x"01010159",
		2692 =>	x"65D5D2D2",
		2693 =>	x"D2D25D59",
		2694 =>	x"01010101",
		2695 =>	x"01010159",
		2696 =>	x"59D3D2D2",
		2697 =>	x"D2D25B59",
		2698 =>	x"01010101",
		2699 =>	x"01010159",
		2700 =>	x"59D6D2D2",
		2701 =>	x"D2D25B59",
		2702 =>	x"01010101",
		2703 =>	x"01010159",
		2704 =>	x"D7D8D2D2",
		2705 =>	x"D2D95D59",
		2706 =>	x"01010101",
		2707 =>	x"01010159",
		2708 =>	x"DAD2D2D2",
		2709 =>	x"D2DB5D59",
		2710 =>	x"01010101",
		2711 =>	x"01015C59",
		2712 =>	x"DCD2D2D2",
		2713 =>	x"D2D25959",
		2714 =>	x"01010101",
		2715 =>	x"01010159",
		2716 =>	x"DDD2D2D2",
		2717 =>	x"D2D25B59",
		2718 =>	x"01010101",
		2719 =>	x"01010159",
		2720 =>	x"59D2D2D2",
		2721 =>	x"D2D26159",
		2722 =>	x"DE010101",
		2723 =>	x"01010159",
		2724 =>	x"DFD2D2D2",
		2725 =>	x"D2E05959",
		2726 =>	x"01010101",
		2727 =>	x"01010159",
		2728 =>	x"DFD3D2D2",
		2729 =>	x"D2E15959",
		2730 =>	x"01010101",
		2731 =>	x"01010159",
		2732 =>	x"59D5D2D2",
		2733 =>	x"D2026159",
		2734 =>	x"DE010101",
		2735 =>	x"01010159",
		2736 =>	x"65D3D2D2",
		2737 =>	x"D2025B59",
		2738 =>	x"01010101",
		2739 =>	x"01010159",
		2740 =>	x"59E2D2D2",
		2741 =>	x"D65F5959",
		2742 =>	x"01010101",
		2743 =>	x"01010101",
		2744 =>	x"59650293",
		2745 =>	x"59595959",
		2746 =>	x"01010101",
		2747 =>	x"01010101",
		2748 =>	x"01595959",
		2749 =>	x"5959E301",
		2750 =>	x"01010101",
		2751 =>	x"01010159", -- IMG_16x16_6intersection
		2752 =>	x"5959E4D2",
		2753 =>	x"D2D2D359",
		2754 =>	x"59010101",
		2755 =>	x"01010159",
		2756 =>	x"5959D5D2",
		2757 =>	x"D2D2D259",
		2758 =>	x"59010101",
		2759 =>	x"0101015C",
		2760 =>	x"5902D2D2",
		2761 =>	x"D2D2D259",
		2762 =>	x"59010101",
		2763 =>	x"01010159",
		2764 =>	x"5902D2D2",
		2765 =>	x"D2D2D259",
		2766 =>	x"59010101",
		2767 =>	x"595959D2",
		2768 =>	x"D2D2D2D2",
		2769 =>	x"D2D2D2D2",
		2770 =>	x"D2595959",
		2771 =>	x"6D59E5D5",
		2772 =>	x"D2D2D2D2",
		2773 =>	x"D2D2D2D3",
		2774 =>	x"D2656502",
		2775 =>	x"D5D5D2D2",
		2776 =>	x"D2D2D2D2",
		2777 =>	x"D2D2D2D2",
		2778 =>	x"D2D5D1D5",
		2779 =>	x"D2D2D2D2",
		2780 =>	x"D2D2D2D2",
		2781 =>	x"D2E6D2D2",
		2782 =>	x"D2E6D2D2",
		2783 =>	x"D2D2D2D2",
		2784 =>	x"D2D2D2D2",
		2785 =>	x"E6D2D2D2",
		2786 =>	x"D2D2D2D2",
		2787 =>	x"D2D2D2D2",
		2788 =>	x"D2D2D2D2",
		2789 =>	x"D2D2D2D2",
		2790 =>	x"D2D2D2D9",
		2791 =>	x"E7D2D2D2",
		2792 =>	x"D2D2D2D2",
		2793 =>	x"D2D2D2D2",
		2794 =>	x"D2D25D61",
		2795 =>	x"59595B5B",
		2796 =>	x"71D2D2D2",
		2797 =>	x"D2D2D271",
		2798 =>	x"5B595959",
		2799 =>	x"59595959",
		2800 =>	x"5902D2D2",
		2801 =>	x"D2D2D259",
		2802 =>	x"59595959",
		2803 =>	x"01010159",
		2804 =>	x"597202D2",
		2805 =>	x"D2D2D259",
		2806 =>	x"01010101",
		2807 =>	x"01010159",
		2808 =>	x"595902D2",
		2809 =>	x"D2D2D259",
		2810 =>	x"59010101",
		2811 =>	x"010101E8",
		2812 =>	x"595902D2",
		2813 =>	x"D2D2D659",
		2814 =>	x"59010101",
		2815 =>	x"09000000", -- IMG_16x16_6middle_horizontal
		2816 =>	x"000A0000",
		2817 =>	x"0B0C0000",
		2818 =>	x"00000D0E",
		2819 =>	x"000A0000",
		2820 =>	x"0F101112",
		2821 =>	x"13141516",
		2822 =>	x"00000000",
		2823 =>	x"00000000",
		2824 =>	x"00000000",
		2825 =>	x"00001718",
		2826 =>	x"191A1B1C",
		2827 =>	x"00001B1B",
		2828 =>	x"1D1E1F20",
		2829 =>	x"00000000",
		2830 =>	x"00000000",
		2831 =>	x"00000000",
		2832 =>	x"00000000",
		2833 =>	x"00000000",
		2834 =>	x"00000000",
		2835 =>	x"00000000",
		2836 =>	x"00000000",
		2837 =>	x"00000000",
		2838 =>	x"00000000",
		2839 =>	x"00000000",
		2840 =>	x"00212223",
		2841 =>	x"24252600",
		2842 =>	x"00000000",
		2843 =>	x"00000000",
		2844 =>	x"00000000",
		2845 =>	x"00000000",
		2846 =>	x"00000000",
		2847 =>	x"00000000",
		2848 =>	x"00000000",
		2849 =>	x"00000000",
		2850 =>	x"00000000",
		2851 =>	x"00000000",
		2852 =>	x"00000000",
		2853 =>	x"00000000",
		2854 =>	x"00000000",
		2855 =>	x"00000000",
		2856 =>	x"00000000",
		2857 =>	x"00000000",
		2858 =>	x"00000000",
		2859 =>	x"00000000",
		2860 =>	x"00000000",
		2861 =>	x"00000000",
		2862 =>	x"00000000",
		2863 =>	x"27272727",
		2864 =>	x"27272727",
		2865 =>	x"54555657",
		2866 =>	x"58000000",
		2867 =>	x"27272727",
		2868 =>	x"27272727",
		2869 =>	x"27272727",
		2870 =>	x"27272727",
		2871 =>	x"27272727",
		2872 =>	x"27272727",
		2873 =>	x"27272727",
		2874 =>	x"27272727",
		2875 =>	x"2C2D2E2F",
		2876 =>	x"301E2A2B",
		2877 =>	x"27272727",
		2878 =>	x"27272727",
		2879 =>	x"01010159", -- IMG_16x16_6middle_vertical
		2880 =>	x"59D2E9E9",
		2881 =>	x"E9E9EA59",
		2882 =>	x"EB010101",
		2883 =>	x"01010101",
		2884 =>	x"59E9E9E9",
		2885 =>	x"E9E9E959",
		2886 =>	x"EB010101",
		2887 =>	x"010101EC",
		2888 =>	x"59E9E9E9",
		2889 =>	x"E9E9E959",
		2890 =>	x"EB010101",
		2891 =>	x"010101EC",
		2892 =>	x"5959E9E9",
		2893 =>	x"E9E9E959",
		2894 =>	x"59010101",
		2895 =>	x"01010159",
		2896 =>	x"59E9E9E9",
		2897 =>	x"E9E95959",
		2898 =>	x"EB010101",
		2899 =>	x"01010159",
		2900 =>	x"59E9E9E9",
		2901 =>	x"E9E9E992",
		2902 =>	x"59010101",
		2903 =>	x"010101EC",
		2904 =>	x"59E9E9E9",
		2905 =>	x"E9E9E992",
		2906 =>	x"59010101",
		2907 =>	x"01010159",
		2908 =>	x"59E9E9E9",
		2909 =>	x"E9E95959",
		2910 =>	x"59010101",
		2911 =>	x"01010159",
		2912 =>	x"59E9E9E9",
		2913 =>	x"E9E9E959",
		2914 =>	x"59010101",
		2915 =>	x"01010159",
		2916 =>	x"59E9E9E9",
		2917 =>	x"E9E9E959",
		2918 =>	x"59010101",
		2919 =>	x"01010159",
		2920 =>	x"9259E9E9",
		2921 =>	x"E9E9E959",
		2922 =>	x"EB010101",
		2923 =>	x"010101EC",
		2924 =>	x"92E9E9E9",
		2925 =>	x"E9E9E959",
		2926 =>	x"EB010101",
		2927 =>	x"010101EC",
		2928 =>	x"59E9E9E9",
		2929 =>	x"E9E9E959",
		2930 =>	x"59010101",
		2931 =>	x"01010101",
		2932 =>	x"59E9E9E9",
		2933 =>	x"E9E95959",
		2934 =>	x"59010101",
		2935 =>	x"01010159",
		2936 =>	x"92E6E9E9",
		2937 =>	x"E9E9E959",
		2938 =>	x"59010101",
		2939 =>	x"01010159",
		2940 =>	x"92D2E9E9",
		2941 =>	x"E9E9E959",
		2942 =>	x"59010101",
		2943 =>	x"01010101", -- IMG_16x16_7end_down
		2944 =>	x"6B593535",
		2945 =>	x"025F5959",
		2946 =>	x"01010101",
		2947 =>	x"01010164",
		2948 =>	x"59653535",
		2949 =>	x"025F5959",
		2950 =>	x"01010101",
		2951 =>	x"01010101",
		2952 =>	x"01653535",
		2953 =>	x"35595901",
		2954 =>	x"01010101",
		2955 =>	x"01010164",
		2956 =>	x"59593535",
		2957 =>	x"355B5901",
		2958 =>	x"01010101",
		2959 =>	x"01010101",
		2960 =>	x"6B593535",
		2961 =>	x"355F5901",
		2962 =>	x"01010101",
		2963 =>	x"01010101",
		2964 =>	x"59653535",
		2965 =>	x"35590101",
		2966 =>	x"01010101",
		2967 =>	x"01010101",
		2968 =>	x"6B653535",
		2969 =>	x"025B5901",
		2970 =>	x"01010101",
		2971 =>	x"01010164",
		2972 =>	x"59593535",
		2973 =>	x"025B5901",
		2974 =>	x"01010101",
		2975 =>	x"01010101",
		2976 =>	x"59593535",
		2977 =>	x"025B0101",
		2978 =>	x"01010101",
		2979 =>	x"01010101",
		2980 =>	x"59353535",
		2981 =>	x"5B595901",
		2982 =>	x"01010101",
		2983 =>	x"01010101",
		2984 =>	x"59593535",
		2985 =>	x"93590101",
		2986 =>	x"01010101",
		2987 =>	x"01010101",
		2988 =>	x"59593535",
		2989 =>	x"355B0101",
		2990 =>	x"01010101",
		2991 =>	x"01010101",
		2992 =>	x"01653535",
		2993 =>	x"35590101",
		2994 =>	x"01010101",
		2995 =>	x"01010101",
		2996 =>	x"59353535",
		2997 =>	x"ED595901",
		2998 =>	x"01010101",
		2999 =>	x"01010101",
		3000 =>	x"01595959",
		3001 =>	x"59590101",
		3002 =>	x"01010101",
		3003 =>	x"01010101",
		3004 =>	x"01010101",
		3005 =>	x"01010101",
		3006 =>	x"01010101",
		3007 =>	x"09000000", -- IMG_16x16_7end_left
		3008 =>	x"000A0000",
		3009 =>	x"0B0C0000",
		3010 =>	x"00000D0E",
		3011 =>	x"000A0000",
		3012 =>	x"0F101112",
		3013 =>	x"13141516",
		3014 =>	x"00000000",
		3015 =>	x"00000000",
		3016 =>	x"00000000",
		3017 =>	x"00001718",
		3018 =>	x"191A1B1C",
		3019 =>	x"00001B1B",
		3020 =>	x"1D1E1F20",
		3021 =>	x"00000000",
		3022 =>	x"00000000",
		3023 =>	x"00000000",
		3024 =>	x"00000000",
		3025 =>	x"00000000",
		3026 =>	x"00000000",
		3027 =>	x"00000000",
		3028 =>	x"00000000",
		3029 =>	x"00000000",
		3030 =>	x"00000000",
		3031 =>	x"00000000",
		3032 =>	x"00212223",
		3033 =>	x"24252600",
		3034 =>	x"00000000",
		3035 =>	x"00000000",
		3036 =>	x"00000000",
		3037 =>	x"00000000",
		3038 =>	x"00000000",
		3039 =>	x"00000000",
		3040 =>	x"00000000",
		3041 =>	x"00000000",
		3042 =>	x"00000000",
		3043 =>	x"00000000",
		3044 =>	x"00000000",
		3045 =>	x"00000000",
		3046 =>	x"00000000",
		3047 =>	x"00000000",
		3048 =>	x"00000000",
		3049 =>	x"00000000",
		3050 =>	x"00000000",
		3051 =>	x"00000000",
		3052 =>	x"00000000",
		3053 =>	x"00000000",
		3054 =>	x"00000000",
		3055 =>	x"27273128",
		3056 =>	x"291E2A2B",
		3057 =>	x"54555657",
		3058 =>	x"58000000",
		3059 =>	x"27272727",
		3060 =>	x"27272727",
		3061 =>	x"27272727",
		3062 =>	x"27272727",
		3063 =>	x"27272727",
		3064 =>	x"27272727",
		3065 =>	x"27272727",
		3066 =>	x"27272727",
		3067 =>	x"2C2D2E2F",
		3068 =>	x"301E2A2B",
		3069 =>	x"27272727",
		3070 =>	x"27272727",
		3071 =>	x"09000000", -- IMG_16x16_7end_right
		3072 =>	x"000A0000",
		3073 =>	x"0B0C0000",
		3074 =>	x"00000D0E",
		3075 =>	x"000A0000",
		3076 =>	x"0F101112",
		3077 =>	x"13141516",
		3078 =>	x"00000000",
		3079 =>	x"00000000",
		3080 =>	x"00000000",
		3081 =>	x"00001718",
		3082 =>	x"191A1B1C",
		3083 =>	x"00001B1B",
		3084 =>	x"1D1E1F20",
		3085 =>	x"00000000",
		3086 =>	x"00000000",
		3087 =>	x"00000000",
		3088 =>	x"00000000",
		3089 =>	x"00000000",
		3090 =>	x"00000000",
		3091 =>	x"00000000",
		3092 =>	x"00000000",
		3093 =>	x"00000000",
		3094 =>	x"00000000",
		3095 =>	x"00000000",
		3096 =>	x"00212223",
		3097 =>	x"24252600",
		3098 =>	x"00000000",
		3099 =>	x"00000000",
		3100 =>	x"00000000",
		3101 =>	x"00000000",
		3102 =>	x"00000000",
		3103 =>	x"00000000",
		3104 =>	x"00000000",
		3105 =>	x"00000000",
		3106 =>	x"00000000",
		3107 =>	x"00000000",
		3108 =>	x"00000000",
		3109 =>	x"00000000",
		3110 =>	x"00000000",
		3111 =>	x"00000000",
		3112 =>	x"00000000",
		3113 =>	x"00000000",
		3114 =>	x"00000000",
		3115 =>	x"00000000",
		3116 =>	x"00000000",
		3117 =>	x"00000000",
		3118 =>	x"00000000",
		3119 =>	x"27273128",
		3120 =>	x"291E2A2B",
		3121 =>	x"54555657",
		3122 =>	x"58000000",
		3123 =>	x"27272727",
		3124 =>	x"27272727",
		3125 =>	x"27272727",
		3126 =>	x"27272727",
		3127 =>	x"27272727",
		3128 =>	x"27272727",
		3129 =>	x"27272727",
		3130 =>	x"27272727",
		3131 =>	x"2C2D2E2F",
		3132 =>	x"301E2A2B",
		3133 =>	x"27272727",
		3134 =>	x"27272727",
		3135 =>	x"09000000", -- IMG_16x16_7end_up
		3136 =>	x"000A0000",
		3137 =>	x"0B0C0000",
		3138 =>	x"00000D0E",
		3139 =>	x"000A0000",
		3140 =>	x"0F101112",
		3141 =>	x"13141516",
		3142 =>	x"00000000",
		3143 =>	x"00000000",
		3144 =>	x"00000000",
		3145 =>	x"00001718",
		3146 =>	x"191A1B1C",
		3147 =>	x"00001B1B",
		3148 =>	x"1D1E1F20",
		3149 =>	x"00000000",
		3150 =>	x"00000000",
		3151 =>	x"00000000",
		3152 =>	x"00000000",
		3153 =>	x"00000000",
		3154 =>	x"00000000",
		3155 =>	x"00000000",
		3156 =>	x"00000000",
		3157 =>	x"00000000",
		3158 =>	x"00000000",
		3159 =>	x"00000000",
		3160 =>	x"00212223",
		3161 =>	x"24252600",
		3162 =>	x"00000000",
		3163 =>	x"00000000",
		3164 =>	x"00000000",
		3165 =>	x"00000000",
		3166 =>	x"00000000",
		3167 =>	x"00000000",
		3168 =>	x"00000000",
		3169 =>	x"00000000",
		3170 =>	x"00000000",
		3171 =>	x"00000000",
		3172 =>	x"00000000",
		3173 =>	x"00000000",
		3174 =>	x"00000000",
		3175 =>	x"00000000",
		3176 =>	x"00000000",
		3177 =>	x"00000000",
		3178 =>	x"00000000",
		3179 =>	x"00000000",
		3180 =>	x"00000000",
		3181 =>	x"00000000",
		3182 =>	x"00000000",
		3183 =>	x"27273128",
		3184 =>	x"291E2A2B",
		3185 =>	x"54555657",
		3186 =>	x"58000000",
		3187 =>	x"27272727",
		3188 =>	x"27272727",
		3189 =>	x"27272727",
		3190 =>	x"27272727",
		3191 =>	x"27272727",
		3192 =>	x"27272727",
		3193 =>	x"27272727",
		3194 =>	x"27272727",
		3195 =>	x"2C2D2E2F",
		3196 =>	x"301E2A2B",
		3197 =>	x"27272727",
		3198 =>	x"27272727",
		3199 =>	x"01010101", -- IMG_16x16_7middle_horizontal
		3200 =>	x"01010101",
		3201 =>	x"01010101",
		3202 =>	x"01010101",
		3203 =>	x"01010101",
		3204 =>	x"01010101",
		3205 =>	x"01010101",
		3206 =>	x"01010101",
		3207 =>	x"01010101",
		3208 =>	x"01010101",
		3209 =>	x"01010101",
		3210 =>	x"01010101",
		3211 =>	x"01010101",
		3212 =>	x"01010101",
		3213 =>	x"01010101",
		3214 =>	x"01010101",
		3215 =>	x"59590159",
		3216 =>	x"59015901",
		3217 =>	x"01010101",
		3218 =>	x"01010101",
		3219 =>	x"59595959",
		3220 =>	x"59595959",
		3221 =>	x"EE595959",
		3222 =>	x"EE59EE59",
		3223 =>	x"EFF0F0F0",
		3224 =>	x"F0F0F0F1",
		3225 =>	x"F2F3F4F0",
		3226 =>	x"F0F0F0F4",
		3227 =>	x"F0F0F0F0",
		3228 =>	x"F0F0F0F0",
		3229 =>	x"F0F0F0F0",
		3230 =>	x"F0F0F0F0",
		3231 =>	x"F0F0F0F0",
		3232 =>	x"F0F0F0F0",
		3233 =>	x"F0F0F0F0",
		3234 =>	x"F0F0F0F0",
		3235 =>	x"F0F0F0F0",
		3236 =>	x"F0F0F0F0",
		3237 =>	x"F0F0F0F0",
		3238 =>	x"F0F0F0F0",
		3239 =>	x"59595959",
		3240 =>	x"59595959",
		3241 =>	x"59F55959",
		3242 =>	x"59595959",
		3243 =>	x"01590159",
		3244 =>	x"01590159",
		3245 =>	x"F6F65959",
		3246 =>	x"01590101",
		3247 =>	x"01010101",
		3248 =>	x"01010101",
		3249 =>	x"01010101",
		3250 =>	x"01010101",
		3251 =>	x"01010101",
		3252 =>	x"01010101",
		3253 =>	x"01010101",
		3254 =>	x"01010101",
		3255 =>	x"01010101",
		3256 =>	x"01010101",
		3257 =>	x"01010101",
		3258 =>	x"01010101",
		3259 =>	x"01010101",
		3260 =>	x"01010101",
		3261 =>	x"01010101",
		3262 =>	x"01010101",
		3263 =>	x"09000000", -- IMG_16x16_7middle_vertical
		3264 =>	x"000A0000",
		3265 =>	x"0B0C0000",
		3266 =>	x"00000D0E",
		3267 =>	x"000A0000",
		3268 =>	x"0F101112",
		3269 =>	x"13141516",
		3270 =>	x"00000000",
		3271 =>	x"00000000",
		3272 =>	x"00000000",
		3273 =>	x"00001718",
		3274 =>	x"191A1B1C",
		3275 =>	x"00001B1B",
		3276 =>	x"1D1E1F20",
		3277 =>	x"00000000",
		3278 =>	x"00000000",
		3279 =>	x"00000000",
		3280 =>	x"00000000",
		3281 =>	x"00000000",
		3282 =>	x"00000000",
		3283 =>	x"00000000",
		3284 =>	x"00000000",
		3285 =>	x"00000000",
		3286 =>	x"00000000",
		3287 =>	x"00000000",
		3288 =>	x"00212223",
		3289 =>	x"24252600",
		3290 =>	x"00000000",
		3291 =>	x"00000000",
		3292 =>	x"00000000",
		3293 =>	x"00000000",
		3294 =>	x"00000000",
		3295 =>	x"00000000",
		3296 =>	x"00000000",
		3297 =>	x"00000000",
		3298 =>	x"00000000",
		3299 =>	x"00000000",
		3300 =>	x"00000000",
		3301 =>	x"00000000",
		3302 =>	x"00000000",
		3303 =>	x"00000000",
		3304 =>	x"00000000",
		3305 =>	x"00000000",
		3306 =>	x"00000000",
		3307 =>	x"00000000",
		3308 =>	x"00000000",
		3309 =>	x"00000000",
		3310 =>	x"00000000",
		3311 =>	x"27272727",
		3312 =>	x"27272727",
		3313 =>	x"54555657",
		3314 =>	x"58000000",
		3315 =>	x"27272727",
		3316 =>	x"27272727",
		3317 =>	x"27272727",
		3318 =>	x"27272727",
		3319 =>	x"27272727",
		3320 =>	x"27272727",
		3321 =>	x"27272727",
		3322 =>	x"27272727",
		3323 =>	x"2C2D2E2F",
		3324 =>	x"301E2A2B",
		3325 =>	x"27272727",
		3326 =>	x"27272727",
		3327 =>	x"F7F7F7F7", -- IMG_16x16_background
		3328 =>	x"F7F7F7F7",
		3329 =>	x"F7F7F7F7",
		3330 =>	x"F7F7F7F7",
		3331 =>	x"F7F7F7F7",
		3332 =>	x"F7F7F7F7",
		3333 =>	x"F7F7F7F7",
		3334 =>	x"F7F7F7F7",
		3335 =>	x"F7F7F7F7",
		3336 =>	x"F7F7F7F7",
		3337 =>	x"F7F7F7F7",
		3338 =>	x"F7F7F7F7",
		3339 =>	x"F7F7F7F7",
		3340 =>	x"F7F7F7F7",
		3341 =>	x"F7F7F7F7",
		3342 =>	x"F7F7F7F7",
		3343 =>	x"F7F7F7F7",
		3344 =>	x"F7F7F7F7",
		3345 =>	x"F7F7F7F7",
		3346 =>	x"F7F7F7F7",
		3347 =>	x"F7F7F7F7",
		3348 =>	x"F7F7F7F7",
		3349 =>	x"F7F7F7F7",
		3350 =>	x"F7F7F7F7",
		3351 =>	x"F7F7F7F7",
		3352 =>	x"F7F7F7F7",
		3353 =>	x"F7F7F7F7",
		3354 =>	x"F7F7F7F7",
		3355 =>	x"F7F7F7F7",
		3356 =>	x"F7F7F7F7",
		3357 =>	x"F7F7F7F7",
		3358 =>	x"F7F7F7F7",
		3359 =>	x"F7F7F7F7",
		3360 =>	x"F7F7F7F7",
		3361 =>	x"F7F7F7F7",
		3362 =>	x"F7F7F7F7",
		3363 =>	x"F7F7F7F7",
		3364 =>	x"F7F7F7F7",
		3365 =>	x"F7F7F7F7",
		3366 =>	x"F7F7F7F7",
		3367 =>	x"F7F7F7F7",
		3368 =>	x"F7F7F7F7",
		3369 =>	x"F7F7F7F7",
		3370 =>	x"F7F7F7F7",
		3371 =>	x"F7F7F7F7",
		3372 =>	x"F7F7F7F7",
		3373 =>	x"F7F7F7F7",
		3374 =>	x"F7F7F7F7",
		3375 =>	x"F7F7F7F7",
		3376 =>	x"F7F7F7F7",
		3377 =>	x"F7F7F7F7",
		3378 =>	x"F7F7F7F7",
		3379 =>	x"F7F7F7F7",
		3380 =>	x"F7F7F7F7",
		3381 =>	x"F7F7F7F7",
		3382 =>	x"F7F7F7F7",
		3383 =>	x"F7F7F7F7",
		3384 =>	x"F7F7F7F7",
		3385 =>	x"F7F7F7F7",
		3386 =>	x"F7F7F7F7",
		3387 =>	x"F7F7F7F7",
		3388 =>	x"F7F7F7F7",
		3389 =>	x"F7F7F7F7",
		3390 =>	x"F7F7F7F7",
		3391 =>	x"01010101", -- IMG_16x16_block
		3392 =>	x"01010101",
		3393 =>	x"01010101",
		3394 =>	x"0101F8F7",
		3395 =>	x"F9F9F9F9",
		3396 =>	x"F9F9F9F9",
		3397 =>	x"F9F9F9F9",
		3398 =>	x"F9F9F8F7",
		3399 =>	x"F9F9F9F9",
		3400 =>	x"F9F9F9F9",
		3401 =>	x"F9F9F9F9",
		3402 =>	x"F9F9F8F7",
		3403 =>	x"F9F9F9F9",
		3404 =>	x"F9F9F9F9",
		3405 =>	x"F9F9F9F9",
		3406 =>	x"F9F9F8F7",
		3407 =>	x"F9F9F9F9",
		3408 =>	x"F9F9F9F9",
		3409 =>	x"F9F9F9F9",
		3410 =>	x"F9F9F8F7",
		3411 =>	x"F9F9F9F9",
		3412 =>	x"F9F9F9F9",
		3413 =>	x"F9F9F9F9",
		3414 =>	x"F9F9F8F7",
		3415 =>	x"F9F9F9F9",
		3416 =>	x"F9F9F9F9",
		3417 =>	x"F9F9F9F9",
		3418 =>	x"F9F9F8F7",
		3419 =>	x"F9F9F9F9",
		3420 =>	x"F9F9F9F9",
		3421 =>	x"F9F9F9F9",
		3422 =>	x"F9F9F8F7",
		3423 =>	x"F9F9F9F9",
		3424 =>	x"F9F9F9F9",
		3425 =>	x"F9F9F9F9",
		3426 =>	x"F9F9F8F7",
		3427 =>	x"F9F9F9F9",
		3428 =>	x"F9F9F9F9",
		3429 =>	x"F9F9F9F9",
		3430 =>	x"F9F9F8F7",
		3431 =>	x"F9F9F9F9",
		3432 =>	x"F9F9F9F9",
		3433 =>	x"F9F9F9F9",
		3434 =>	x"F9F9F8F7",
		3435 =>	x"F9F9F9F9",
		3436 =>	x"F9F9F9F9",
		3437 =>	x"F9F9F9F9",
		3438 =>	x"F9F9F8F7",
		3439 =>	x"F9F9F9F9",
		3440 =>	x"F9F9F9F9",
		3441 =>	x"F9F9F9F9",
		3442 =>	x"F9F9F8F7",
		3443 =>	x"F9F9F9F9",
		3444 =>	x"F9F9F9F9",
		3445 =>	x"F9F9F9F9",
		3446 =>	x"F9F9F8F7",
		3447 =>	x"F8F8F8F8",
		3448 =>	x"F8F8F8F8",
		3449 =>	x"F8F8F8F8",
		3450 =>	x"F8F9F8F7",
		3451 =>	x"F8F8F8F8",
		3452 =>	x"F8F8F8F8",
		3453 =>	x"F8F8F8F8",
		3454 =>	x"F8F8F8F7",
		3455 =>	x"F7F7F7F7", -- IMG_16x16_bomb
		3456 =>	x"F7F7F7F7",
		3457 =>	x"F7F7F7F7",
		3458 =>	x"F7F7F7F7",
		3459 =>	x"F7F7F7F7",
		3460 =>	x"F7F7F7F7",
		3461 =>	x"F7010101",
		3462 =>	x"F701F701",
		3463 =>	x"F7F7F7F7",
		3464 =>	x"F7F8F8F8",
		3465 =>	x"0101F8F8",
		3466 =>	x"F7F7F7F7",
		3467 =>	x"F7F7F7F8",
		3468 =>	x"F8F8F8F8",
		3469 =>	x"01F8F8F8",
		3470 =>	x"F8F701F7",
		3471 =>	x"F7F7F8F8",
		3472 =>	x"0101F8F8",
		3473 =>	x"01F8F8F8",
		3474 =>	x"F8F8F7F7",
		3475 =>	x"F7F8F801",
		3476 =>	x"01F8F8F8",
		3477 =>	x"F8F8F8F8",
		3478 =>	x"F8F8F8F7",
		3479 =>	x"F7F8F801",
		3480 =>	x"01F8F8F8",
		3481 =>	x"F8F8F8F8",
		3482 =>	x"F8F8F8F7",
		3483 =>	x"F8F80101",
		3484 =>	x"F8F8F8F8",
		3485 =>	x"F8F8F8F8",
		3486 =>	x"F8F8F8F8",
		3487 =>	x"F8F80101",
		3488 =>	x"F8F8F8F8",
		3489 =>	x"F8F8F8F8",
		3490 =>	x"F8F8F8F8",
		3491 =>	x"F8F8F8F8",
		3492 =>	x"F8F8F8F8",
		3493 =>	x"F8F8F8F8",
		3494 =>	x"F8F8F8F8",
		3495 =>	x"F8F8F8F8",
		3496 =>	x"F8F8F8F8",
		3497 =>	x"F8F8F8F8",
		3498 =>	x"F8F8F8F8",
		3499 =>	x"F8F8F8F8",
		3500 =>	x"F8F8F8F8",
		3501 =>	x"F8F8F8F8",
		3502 =>	x"F8F8F8F8",
		3503 =>	x"F7F8F8F8",
		3504 =>	x"F8F8F8F8",
		3505 =>	x"F8F8F8F8",
		3506 =>	x"F8F8F8F7",
		3507 =>	x"F7F8F8F8",
		3508 =>	x"F8F8F8F8",
		3509 =>	x"F8F8F8F8",
		3510 =>	x"F8F8F8F7",
		3511 =>	x"F7F7F8F8",
		3512 =>	x"F8F8F8F8",
		3513 =>	x"F8F8F8F8",
		3514 =>	x"F8F8F7F7",
		3515 =>	x"F7F7F7F8",
		3516 =>	x"F8F8F8F8",
		3517 =>	x"F8F8F8F8",
		3518 =>	x"F8F7F7F7",
		3519 =>	x"F7F7F7F7", -- IMG_16x16_bomberman
		3520 =>	x"F7010101",
		3521 =>	x"010101F7",
		3522 =>	x"F7F7F7F7",
		3523 =>	x"F7F7F7F7",
		3524 =>	x"01010101",
		3525 =>	x"01010101",
		3526 =>	x"F7F7F7F7",
		3527 =>	x"F7F7F7F7",
		3528 =>	x"01FAF7FA",
		3529 =>	x"FAF7FA01",
		3530 =>	x"F7F7F7F7",
		3531 =>	x"F7F7F7F7",
		3532 =>	x"01FAF7FA",
		3533 =>	x"FAF7FA01",
		3534 =>	x"F7F7F7F7",
		3535 =>	x"F7F7F7F7",
		3536 =>	x"01010101",
		3537 =>	x"01010101",
		3538 =>	x"F7F7F7F7",
		3539 =>	x"F7F7F7F7",
		3540 =>	x"F7010101",
		3541 =>	x"010101F7",
		3542 =>	x"F7F7F7F7",
		3543 =>	x"F7F7F7F7",
		3544 =>	x"F7F7FBFB",
		3545 =>	x"FBFBF7F7",
		3546 =>	x"F7F7F7F7",
		3547 =>	x"F7F7F7F7",
		3548 =>	x"0101FBFB",
		3549 =>	x"FBFB0101",
		3550 =>	x"F7F7F7F7",
		3551 =>	x"F7F7F701",
		3552 =>	x"01FBFBFB",
		3553 =>	x"FBFBFB01",
		3554 =>	x"01F7F7F7",
		3555 =>	x"F7F7FAFA",
		3556 =>	x"01FBFBFB",
		3557 =>	x"FBFBFB01",
		3558 =>	x"FAFAF7F7",
		3559 =>	x"F7F7FAFA",
		3560 =>	x"F7FBFBFB",
		3561 =>	x"FBFBFBF7",
		3562 =>	x"FAFAF7F7",
		3563 =>	x"F7F7F7F7",
		3564 =>	x"F7FBFBFB",
		3565 =>	x"FBFBFBF7",
		3566 =>	x"F7F7F7F7",
		3567 =>	x"F7F7F7F7",
		3568 =>	x"F70101FB",
		3569 =>	x"FB0101F7",
		3570 =>	x"F7F7F7F7",
		3571 =>	x"F7F7F7F7",
		3572 =>	x"F70101F7",
		3573 =>	x"F70101F7",
		3574 =>	x"F7F7F7F7",
		3575 =>	x"F7F7F7F7",
		3576 =>	x"F7FAFAF7",
		3577 =>	x"F7FAFAF7",
		3578 =>	x"F7F7F7F7",
		3579 =>	x"F7F7F7F7",
		3580 =>	x"F7FAFAF7",
		3581 =>	x"F7FAFAF7",
		3582 =>	x"F7F7F7F7",
		3583 =>	x"F7F7F7F7", -- IMG_16x16_bomberman_bomb
		3584 =>	x"F7010101",
		3585 =>	x"010101F7",
		3586 =>	x"F7F7F7F7",
		3587 =>	x"F7F7F7F7",
		3588 =>	x"01010101",
		3589 =>	x"01010101",
		3590 =>	x"F7F7F7F7",
		3591 =>	x"F7F7F7F7",
		3592 =>	x"01FAF7FA",
		3593 =>	x"FAF7FA01",
		3594 =>	x"F7F7F7F7",
		3595 =>	x"F7F7F700",
		3596 =>	x"01FAF7FA",
		3597 =>	x"FAF7FA01",
		3598 =>	x"00F7F7F7",
		3599 =>	x"F7F70000",
		3600 =>	x"01010101",
		3601 =>	x"01010101",
		3602 =>	x"0000F7F7",
		3603 =>	x"F7000000",
		3604 =>	x"00010101",
		3605 =>	x"01010100",
		3606 =>	x"000000F7",
		3607 =>	x"F7000000",
		3608 =>	x"0000FBFB",
		3609 =>	x"FBFB0000",
		3610 =>	x"000000F7",
		3611 =>	x"00000000",
		3612 =>	x"0101FBFB",
		3613 =>	x"FBFB0101",
		3614 =>	x"00000000",
		3615 =>	x"00000001",
		3616 =>	x"01FBFBFB",
		3617 =>	x"FBFBFB01",
		3618 =>	x"01000000",
		3619 =>	x"0000FAFA",
		3620 =>	x"01FBFBFB",
		3621 =>	x"FBFBFB01",
		3622 =>	x"FAFA0000",
		3623 =>	x"0000FAFA",
		3624 =>	x"00FBFBFB",
		3625 =>	x"FBFBFB00",
		3626 =>	x"FAFA0000",
		3627 =>	x"00000000",
		3628 =>	x"00FBFBFB",
		3629 =>	x"FBFBFB00",
		3630 =>	x"00000000",
		3631 =>	x"F7000000",
		3632 =>	x"000101FB",
		3633 =>	x"FB010100",
		3634 =>	x"000000F7",
		3635 =>	x"F7000000",
		3636 =>	x"00010100",
		3637 =>	x"00010100",
		3638 =>	x"000000F7",
		3639 =>	x"F7F70000",
		3640 =>	x"00FAFA00",
		3641 =>	x"00FAFA00",
		3642 =>	x"0000F7F7",
		3643 =>	x"F7F7F700",
		3644 =>	x"00FAFA00",
		3645 =>	x"00FAFA00",
		3646 =>	x"00F7F7F7",
		3647 =>	x"F8F8F8F8", -- IMG_16x16_brick
		3648 =>	x"F8F8F8F8",
		3649 =>	x"F8F8F8F8",
		3650 =>	x"F8F8F8F8",
		3651 =>	x"F8010101",
		3652 =>	x"01010101",
		3653 =>	x"01010101",
		3654 =>	x"010101F8",
		3655 =>	x"01F9F9F9",
		3656 =>	x"F9F9F9F9",
		3657 =>	x"F9F9F9F9",
		3658 =>	x"F9F9F9F8",
		3659 =>	x"01F9F9F9",
		3660 =>	x"F9F9F9F9",
		3661 =>	x"F9F9F9F9",
		3662 =>	x"F9F9F9F8",
		3663 =>	x"01F9F9F9",
		3664 =>	x"F9F9F9F9",
		3665 =>	x"F9F9F9F9",
		3666 =>	x"F9F9F9F8",
		3667 =>	x"F8F8F8F8",
		3668 =>	x"F8F8F8F8",
		3669 =>	x"F8F8F8F8",
		3670 =>	x"F8F8F8F8",
		3671 =>	x"01010101",
		3672 =>	x"01F8F801",
		3673 =>	x"01010101",
		3674 =>	x"01010101",
		3675 =>	x"F9F9F9F9",
		3676 =>	x"F9F801F9",
		3677 =>	x"F9F9F9F9",
		3678 =>	x"F9F9F9F9",
		3679 =>	x"F9F9F9F9",
		3680 =>	x"F9F801F9",
		3681 =>	x"F9F9F9F9",
		3682 =>	x"F9F9F9F9",
		3683 =>	x"F9F9F9F9",
		3684 =>	x"F9F801F9",
		3685 =>	x"F9F9F9F9",
		3686 =>	x"F9F9F9F9",
		3687 =>	x"F8F8F8F8",
		3688 =>	x"F8F8F8F8",
		3689 =>	x"F8F8F8F8",
		3690 =>	x"F8F8F8F8",
		3691 =>	x"01010101",
		3692 =>	x"01010101",
		3693 =>	x"01F8F801",
		3694 =>	x"01010101",
		3695 =>	x"F9F9F9F9",
		3696 =>	x"F9F9F9F9",
		3697 =>	x"F9F801F9",
		3698 =>	x"F9F9F9F9",
		3699 =>	x"F9F9F9F9",
		3700 =>	x"F9F9F9F9",
		3701 =>	x"F9F801F9",
		3702 =>	x"F9F9F9F9",
		3703 =>	x"F9F9F9F9",
		3704 =>	x"F9F9F9F9",
		3705 =>	x"F9F801F9",
		3706 =>	x"F9F9F9F9",
		3707 =>	x"F8F8F8F8",
		3708 =>	x"F8F8F8F8",
		3709 =>	x"F8F8F8F8",
		3710 =>	x"F8F8F8F8",
		3711 =>	x"F8FCFCFC", -- IMG_16x16_door
		3712 =>	x"FCFCF8FC",
		3713 =>	x"FCFCFCFC",
		3714 =>	x"F8F8F7F7",
		3715 =>	x"FCFCFDFD",
		3716 =>	x"FDFCF8FC",
		3717 =>	x"FDFDFDFC",
		3718 =>	x"FCF8F7F7",
		3719 =>	x"FCFDFDFC",
		3720 =>	x"FDFCF8FC",
		3721 =>	x"FDFCFDFD",
		3722 =>	x"FCFCF7F7",
		3723 =>	x"FCFDFDFD",
		3724 =>	x"FDFCF8FC",
		3725 =>	x"FDFDFDFD",
		3726 =>	x"FCFCF7F7",
		3727 =>	x"FCFDFDFD",
		3728 =>	x"FDFCF8FC",
		3729 =>	x"FDFDFDFD",
		3730 =>	x"FCF8F7F7",
		3731 =>	x"FCFDFDF8",
		3732 =>	x"FDFCF8FC",
		3733 =>	x"FDF8FDFD",
		3734 =>	x"FCF8F7F7",
		3735 =>	x"FCFDFCF8",
		3736 =>	x"FCFCFCFC",
		3737 =>	x"FCF8FCFD",
		3738 =>	x"FCF8F7F7",
		3739 =>	x"FCFDFCF8",
		3740 =>	x"FCFCFCFC",
		3741 =>	x"FCF8FCFD",
		3742 =>	x"FCF8F7F7",
		3743 =>	x"FCFDFDF8",
		3744 =>	x"FDFCF8FC",
		3745 =>	x"FDF8FDFD",
		3746 =>	x"FCF8F7F7",
		3747 =>	x"FCFDFDFD",
		3748 =>	x"FDFCF8FC",
		3749 =>	x"FDFDFDFD",
		3750 =>	x"FCF8F7F7",
		3751 =>	x"FCFDFDFD",
		3752 =>	x"FDFCF8FC",
		3753 =>	x"FDFDFDFD",
		3754 =>	x"FCFCF7F7",
		3755 =>	x"FCFDFDFC",
		3756 =>	x"FDFCF8FC",
		3757 =>	x"FDFCFDFD",
		3758 =>	x"FCFCF7F7",
		3759 =>	x"FCFCFDFD",
		3760 =>	x"FDFCF8FC",
		3761 =>	x"FDFDFDFC",
		3762 =>	x"FCF8F7F7",
		3763 =>	x"F8FCFCFC",
		3764 =>	x"FCFCF8FC",
		3765 =>	x"FCFCFCFC",
		3766 =>	x"F8F8F7F7",
		3767 =>	x"F7F7F7F7",
		3768 =>	x"F7F7F7F7",
		3769 =>	x"F7F7F7F7",
		3770 =>	x"F7F7F7F7",
		3771 =>	x"F7F7F7F7",
		3772 =>	x"F7F7F7F7",
		3773 =>	x"F7F7F7F7",
		3774 =>	x"F7F7F7F7",
		3775 =>	x"F7F7F7F7", -- IMG_16x16_enemy
		3776 =>	x"F7F7F7F7",
		3777 =>	x"F7F7F7F7",
		3778 =>	x"F7F7F7F7",
		3779 =>	x"F7F7F7F7",
		3780 =>	x"F7F7F7F7",
		3781 =>	x"F7F7F7F7",
		3782 =>	x"F7F7F7F7",
		3783 =>	x"F7F7F7F7",
		3784 =>	x"F8F8F8F8",
		3785 =>	x"F8F8F8F8",
		3786 =>	x"F7F7F7F7",
		3787 =>	x"F7F7F8F8",
		3788 =>	x"F8FAFAFA",
		3789 =>	x"FAFAFAF8",
		3790 =>	x"F8F8F7F7",
		3791 =>	x"F7F8F8FA",
		3792 =>	x"FAFAFAFA",
		3793 =>	x"FAFAFAFA",
		3794 =>	x"FAF8F8F7",
		3795 =>	x"F8F8FAFA",
		3796 =>	x"FAFAFAFA",
		3797 =>	x"FAFAFAFA",
		3798 =>	x"FAFAF8F8",
		3799 =>	x"F8FAFAFA",
		3800 =>	x"FA0101FA",
		3801 =>	x"FA0101FA",
		3802 =>	x"FAFAFAF8",
		3803 =>	x"F8FAFAFA",
		3804 =>	x"FAF801FA",
		3805 =>	x"FAF801FA",
		3806 =>	x"FAFAFAF8",
		3807 =>	x"F8FAFAFA",
		3808 =>	x"FAF801FA",
		3809 =>	x"FAF801FA",
		3810 =>	x"FAFAFAF8",
		3811 =>	x"F8F8FAFA",
		3812 =>	x"FAFAFAFA",
		3813 =>	x"FAFAFAFA",
		3814 =>	x"FAFAF8F8",
		3815 =>	x"F7F8FAFA",
		3816 =>	x"FAFAFAFA",
		3817 =>	x"FAFAFAFA",
		3818 =>	x"FAFAF8F7",
		3819 =>	x"F7F8F8FA",
		3820 =>	x"FAFAFAF8",
		3821 =>	x"F8FAFAFA",
		3822 =>	x"FAF8F8F7",
		3823 =>	x"F7F7F8F8",
		3824 =>	x"F8FAFAFA",
		3825 =>	x"FAFAFAF8",
		3826 =>	x"F8F8F7F7",
		3827 =>	x"F7F7F7F7",
		3828 =>	x"F8F8F8FA",
		3829 =>	x"FAF8F8F8",
		3830 =>	x"F7F7F7F7",
		3831 =>	x"F7F7F7F7",
		3832 =>	x"F7F7F801",
		3833 =>	x"01F8F7F7",
		3834 =>	x"F7F7F7F7",
		3835 =>	x"F7F7F7F7",
		3836 =>	x"F7F7F8F8",
		3837 =>	x"F8F8F7F7",
		3838 =>	x"F7F7F7F7",
		3839 =>	x"59595959", -- IMG_16x16_plus_bomb
		3840 =>	x"59595959",
		3841 =>	x"59595959",
		3842 =>	x"59595959",
		3843 =>	x"59808080",
		3844 =>	x"80808080",
		3845 =>	x"80010101",
		3846 =>	x"80808059",
		3847 =>	x"59808080",
		3848 =>	x"80F8F8F8",
		3849 =>	x"0101F8F8",
		3850 =>	x"80808059",
		3851 =>	x"598080F8",
		3852 =>	x"F8F8F8F8",
		3853 =>	x"01F8F8F8",
		3854 =>	x"F8808059",
		3855 =>	x"5980F8F8",
		3856 =>	x"0101F8F8",
		3857 =>	x"01F8F8F8",
		3858 =>	x"F8F88059",
		3859 =>	x"59F8F801",
		3860 =>	x"01F8F8F8",
		3861 =>	x"F8F8F8F8",
		3862 =>	x"F8F8F859",
		3863 =>	x"59F8F801",
		3864 =>	x"01F8F8F8",
		3865 =>	x"F8F8F8F8",
		3866 =>	x"F8F8F859",
		3867 =>	x"59F80101",
		3868 =>	x"F8F8F8F8",
		3869 =>	x"F8F8F8F8",
		3870 =>	x"F8F8F859",
		3871 =>	x"59F80101",
		3872 =>	x"F8F8F8F8",
		3873 =>	x"F8F8F8F8",
		3874 =>	x"F8F8F859",
		3875 =>	x"59F8F8F8",
		3876 =>	x"F8F8F8F8",
		3877 =>	x"F8F8F8F8",
		3878 =>	x"F8F8F859",
		3879 =>	x"59F8F8F8",
		3880 =>	x"F8F8F8F8",
		3881 =>	x"F8F8F8F8",
		3882 =>	x"F8F8F859",
		3883 =>	x"59F8F8F8",
		3884 =>	x"F8F8F8F8",
		3885 =>	x"F8F8F8F8",
		3886 =>	x"F8F8F859",
		3887 =>	x"59F8F8F8",
		3888 =>	x"F8F8F8F8",
		3889 =>	x"F8F8F8F8",
		3890 =>	x"F8F8F859",
		3891 =>	x"59F8F8F8",
		3892 =>	x"F8F8F8F8",
		3893 =>	x"F8F8F8F8",
		3894 =>	x"F8F8F859",
		3895 =>	x"5980F8F8",
		3896 =>	x"F8F8F8F8",
		3897 =>	x"F8F8F8F8",
		3898 =>	x"F8F88059",
		3899 =>	x"59595959",
		3900 =>	x"59595959",
		3901 =>	x"59595959",
		3902 =>	x"59595959",
		3903 =>	x"FEFEFEFE", -- IMG_16x16_plus_explosion
		3904 =>	x"FEFEFEFE",
		3905 =>	x"FEFEFEFE",
		3906 =>	x"FEFEFEFE",
		3907 =>	x"FE808080",
		3908 =>	x"80808080",
		3909 =>	x"80808080",
		3910 =>	x"808080FE",
		3911 =>	x"FE808080",
		3912 =>	x"80808059",
		3913 =>	x"59808080",
		3914 =>	x"808080FE",
		3915 =>	x"FE808080",
		3916 =>	x"80808059",
		3917 =>	x"59808080",
		3918 =>	x"808080FE",
		3919 =>	x"FE808080",
		3920 =>	x"80805993",
		3921 =>	x"93598080",
		3922 =>	x"808080FE",
		3923 =>	x"FE808080",
		3924 =>	x"80595993",
		3925 =>	x"93595980",
		3926 =>	x"808080FE",
		3927 =>	x"FE808080",
		3928 =>	x"59599380",
		3929 =>	x"80935959",
		3930 =>	x"808080FE",
		3931 =>	x"FE805959",
		3932 =>	x"93938080",
		3933 =>	x"80809393",
		3934 =>	x"595980FE",
		3935 =>	x"FE805959",
		3936 =>	x"93938080",
		3937 =>	x"80809393",
		3938 =>	x"595980FE",
		3939 =>	x"FE808080",
		3940 =>	x"59599380",
		3941 =>	x"80935959",
		3942 =>	x"808080FE",
		3943 =>	x"FE808080",
		3944 =>	x"80595993",
		3945 =>	x"93595980",
		3946 =>	x"808080FE",
		3947 =>	x"FE808080",
		3948 =>	x"80805993",
		3949 =>	x"93598080",
		3950 =>	x"808080FE",
		3951 =>	x"FE808080",
		3952 =>	x"80808059",
		3953 =>	x"59808080",
		3954 =>	x"808080FE",
		3955 =>	x"FE808080",
		3956 =>	x"80808059",
		3957 =>	x"59808080",
		3958 =>	x"808080FE",
		3959 =>	x"FE808080",
		3960 =>	x"80808080",
		3961 =>	x"80808080",
		3962 =>	x"808080FE",
		3963 =>	x"FEFEFEFE",
		3964 =>	x"FEFEFEFE",
		3965 =>	x"FEFEFEFE",
		3966 =>	x"FEFEFEFE",


--			***** MAP *****


		3967 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3968 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3969 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3970 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3971 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3972 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3973 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3974 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3975 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3976 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3977 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3978 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3979 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3980 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3981 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3982 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3983 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3984 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3985 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3986 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3987 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3988 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3989 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3990 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3991 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3992 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3993 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3994 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3995 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3996 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3997 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3998 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3999 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4000 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4001 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4002 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4003 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4004 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4005 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4006 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4007 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4008 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4009 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4010 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4011 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4012 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4013 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4014 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4015 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4016 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4017 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4018 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4019 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4020 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4021 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4022 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4023 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4024 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4025 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4026 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4027 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4028 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4029 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4030 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4031 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4032 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4033 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4034 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4035 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4036 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4037 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4038 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4039 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4040 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4041 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4042 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4043 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4044 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4045 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4046 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4047 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4048 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4049 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4050 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4051 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4052 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4053 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4054 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4055 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4056 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4057 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4058 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4059 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4060 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4061 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4062 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4063 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4064 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4065 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4066 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4067 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4068 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4069 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4070 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4071 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4072 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4073 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4074 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4075 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4076 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4077 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4078 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4079 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4080 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4081 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4082 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4083 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4084 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4085 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4086 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4087 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4088 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4089 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4090 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4091 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4092 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4093 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4094 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4095 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4096 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4097 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4098 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4099 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4100 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4101 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4102 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4103 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4104 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4105 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4106 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4107 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4108 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4109 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4110 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4111 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4112 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4113 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4114 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4115 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4116 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4117 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4118 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4119 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4120 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4121 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4122 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4123 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4124 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4125 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4126 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4127 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4128 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4129 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4130 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4131 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4132 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4133 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4134 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4135 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4136 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4137 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4138 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4139 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4140 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4141 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4142 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4143 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4144 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4145 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4146 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4147 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4148 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4149 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4150 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4151 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4152 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4153 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4154 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4155 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4156 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4157 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4158 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4159 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4160 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4161 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4162 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4163 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4164 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4165 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4166 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4167 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4168 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4169 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4170 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4171 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4172 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4173 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4174 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4175 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4176 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4177 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4178 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4179 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4180 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4181 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4182 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4183 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4184 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4185 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4186 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4187 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4188 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4189 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4190 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4191 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4192 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4193 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4194 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4195 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4196 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4197 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4198 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4199 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4200 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4201 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4202 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4203 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4204 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4205 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4206 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4207 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4208 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4209 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4210 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4211 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4212 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4213 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4214 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4215 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4216 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4217 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4218 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4219 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4220 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4221 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4222 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4223 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4224 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4225 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4226 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4227 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4228 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4229 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4230 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4231 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4232 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4233 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4234 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4235 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4236 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4237 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4238 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4239 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4240 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4241 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4242 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4243 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4244 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4245 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4246 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4247 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4248 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4249 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4250 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4251 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4252 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4253 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4254 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4255 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4256 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4257 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4258 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4259 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4260 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4261 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4262 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4263 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4264 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4265 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4266 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4267 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4268 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4269 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4270 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4271 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4272 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4273 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4274 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4275 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4276 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4277 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4278 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4279 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4280 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4281 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4282 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4283 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4284 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4285 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4286 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4287 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4288 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4289 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4290 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4291 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4292 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4293 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4294 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4295 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4296 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4297 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4298 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4299 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4300 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4301 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4302 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4303 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4304 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4305 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4306 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4307 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4308 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4309 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4310 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4311 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4312 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4313 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4314 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4315 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4316 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4317 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4318 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4319 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4320 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4321 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4322 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4323 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4324 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4325 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4326 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4327 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4328 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4329 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4330 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4331 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4332 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4333 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4334 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4335 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4336 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4337 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4338 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4339 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4340 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4341 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4342 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4343 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4344 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4345 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4346 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4347 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4348 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4349 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4350 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4351 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4352 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4353 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4354 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4355 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4356 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4357 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4358 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4359 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4360 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4361 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4362 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4363 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4364 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4365 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4366 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4367 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4368 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4369 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4370 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4371 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4372 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4373 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4374 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4375 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4376 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4377 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4378 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4379 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4380 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4381 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4382 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4383 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4384 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4385 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4386 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4387 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4388 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4389 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4390 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4391 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4392 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4393 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4394 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4395 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4396 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4397 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4398 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4399 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4400 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4401 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4402 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4403 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4404 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4405 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4406 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4407 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4408 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4409 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4410 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4411 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4412 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4413 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4414 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4415 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4416 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4417 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4418 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4419 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4420 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4421 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4422 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4423 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4424 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4425 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4426 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4427 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4428 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4429 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4430 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4431 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4432 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4433 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4434 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4435 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4436 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4437 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4438 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4439 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4440 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4441 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4442 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4443 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4444 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4445 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4446 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4447 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4448 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4449 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4450 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4451 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4452 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4453 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4454 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4455 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4456 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4457 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4458 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4459 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4460 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4461 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4462 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4463 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4464 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4465 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4466 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4467 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4468 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4469 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4470 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4471 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4472 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4473 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4474 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4475 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4476 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4477 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4478 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4479 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4480 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4481 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4482 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4483 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4484 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4485 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4486 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4487 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4488 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4489 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4490 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4491 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4492 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4493 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4494 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4495 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4496 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4497 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4498 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4499 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4500 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4501 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4502 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4503 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4504 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4505 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4506 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4507 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4508 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4509 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4510 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4511 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4512 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4513 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4514 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4515 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4516 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4517 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4518 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4519 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4520 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4521 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4522 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4523 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4524 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4525 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4526 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4527 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4528 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4529 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4530 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4531 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4532 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4533 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4534 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4535 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4536 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4537 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4538 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4539 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4540 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4541 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4542 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4543 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4544 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4545 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4546 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4547 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4548 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4549 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4550 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4551 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4552 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4553 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4554 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4555 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4556 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4557 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4558 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4559 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4560 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4561 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4562 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4563 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4564 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4565 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4566 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4567 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4568 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4569 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4570 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4571 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4572 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4573 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4574 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4575 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4576 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4577 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4578 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4579 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4580 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4581 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4582 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4583 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4584 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4585 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4586 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4587 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4588 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4589 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4590 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4591 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4592 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4593 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4594 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4595 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4596 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4597 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4598 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4599 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4600 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4601 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4602 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4603 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4604 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4605 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4606 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4607 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4608 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4609 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4610 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4611 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4612 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4613 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4614 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4615 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4616 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4617 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4618 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4619 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4620 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4621 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4622 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4623 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4624 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4625 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4626 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4627 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4628 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4629 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4630 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4631 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4632 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4633 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4634 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4635 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4636 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4637 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4638 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4639 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4640 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4641 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4642 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4643 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4644 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4645 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4646 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4647 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4648 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4649 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4650 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4651 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4652 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4653 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4654 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4655 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4656 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4657 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4658 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4659 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4660 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4661 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4662 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4663 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4664 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4665 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4666 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4667 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4668 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4669 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4670 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4671 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4672 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4673 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4674 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4675 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4676 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4677 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4678 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4679 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4680 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4681 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4682 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4683 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4684 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4685 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4686 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4687 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4688 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4689 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4690 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4691 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4692 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4693 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4694 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4695 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4696 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4697 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4698 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4699 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4700 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4701 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4702 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4703 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4704 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4705 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4706 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4707 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4708 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4709 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4710 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4711 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4712 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4713 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4714 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4715 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4716 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4717 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4718 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4719 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4720 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4721 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4722 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4723 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4724 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4725 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4726 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4727 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4728 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4729 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4730 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4731 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4732 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4733 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4734 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4735 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4736 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4737 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4738 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4739 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4740 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4741 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4742 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4743 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4744 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4745 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4746 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4747 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4748 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4749 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4750 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4751 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4752 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4753 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4754 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4755 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4756 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4757 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4758 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4759 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4760 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4761 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4762 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4763 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4764 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4765 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4766 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4767 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4768 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4769 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4770 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4771 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4772 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4773 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4774 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4775 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4776 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4777 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4778 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4779 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4780 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4781 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4782 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4783 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4784 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4785 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4786 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4787 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4788 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4789 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4790 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4791 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4792 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4793 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4794 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4795 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4796 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4797 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4798 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4799 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4800 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4801 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4802 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4803 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4804 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4805 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4806 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4807 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4808 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4809 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4810 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4811 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4812 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4813 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4814 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4815 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4816 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4817 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4818 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4819 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4820 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4821 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4822 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4823 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4824 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4825 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4826 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4827 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4828 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4829 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4830 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4831 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4832 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4833 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4834 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4835 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4836 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4837 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4838 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4839 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4840 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4841 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4842 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4843 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4844 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4845 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4846 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4847 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4848 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4849 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4850 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4851 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4852 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4853 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4854 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4855 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4856 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4857 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4858 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4859 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4860 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4861 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4862 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4863 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4864 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4865 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4866 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4867 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4868 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4869 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4870 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4871 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4872 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4873 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4874 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4875 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4876 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4877 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4878 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4879 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4880 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4881 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4882 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4883 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4884 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4885 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4886 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4887 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4888 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4889 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4890 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4891 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4892 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4893 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4894 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4895 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4896 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4897 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4898 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4899 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4900 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4901 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4902 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4903 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4904 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4905 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4906 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4907 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4908 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4909 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4910 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4911 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4912 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4913 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4914 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4915 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4916 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4917 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4918 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4919 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4920 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4921 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4922 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4923 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4924 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4925 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4926 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4927 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4928 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4929 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4930 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4931 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4932 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4933 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4934 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4935 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4936 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4937 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4938 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4939 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4940 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4941 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4942 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4943 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4944 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4945 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4946 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4947 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4948 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4949 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4950 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4951 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4952 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4953 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4954 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4955 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4956 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4957 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4958 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4959 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4960 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4961 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4962 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4963 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4964 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4965 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4966 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4967 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4968 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4969 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4970 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4971 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4972 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4973 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4974 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4975 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4976 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4977 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4978 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4979 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4980 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4981 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4982 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4983 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4984 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4985 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4986 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4987 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4988 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4989 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4990 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4991 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4992 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4993 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4994 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4995 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4996 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4997 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4998 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4999 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5000 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5001 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5002 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5003 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5004 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5005 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5006 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5007 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5008 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5009 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5010 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5011 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5012 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5013 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5014 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5015 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5016 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5017 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5018 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5019 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5020 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5021 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5022 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5023 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5024 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5025 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5026 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5027 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5028 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5029 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5030 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5031 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5032 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5033 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5034 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5035 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5036 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5037 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5038 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5039 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5040 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5041 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5042 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5043 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5044 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5045 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5046 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5047 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5048 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5049 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5050 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5051 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5052 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5053 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5054 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5055 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5056 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5057 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5058 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5059 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5060 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5061 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5062 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5063 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5064 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5065 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5066 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5067 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5068 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5069 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5070 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5071 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5072 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5073 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5074 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5075 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5076 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5077 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5078 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5079 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5080 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5081 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5082 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5083 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5084 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5085 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5086 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5087 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5088 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5089 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5090 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5091 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5092 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5093 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5094 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5095 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5096 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5097 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5098 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5099 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5100 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5101 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5102 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5103 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5104 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5105 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5106 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5107 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5108 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5109 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5110 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5111 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5112 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5113 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5114 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5115 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5116 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5117 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5118 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5119 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5120 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5121 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5122 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5123 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5124 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5125 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5126 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5127 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5128 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5129 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5130 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5131 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5132 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5133 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5134 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5135 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5136 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5137 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5138 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5139 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5140 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5141 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5142 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5143 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5144 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5145 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5146 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5147 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5148 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5149 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5150 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5151 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5152 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5153 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5154 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5155 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5156 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5157 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5158 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5159 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5160 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5161 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5162 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5163 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5164 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5165 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5166 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
			0 =>	x"00000000", -- R: 0 G: 0 B: 0
		1 =>	x"00FFFFFF", -- R: 255 G: 255 B: 255
		2 =>	x"00004DFF", -- R: 255 G: 77 B: 0
		3 =>	x"0044B3FF", -- R: 255 G: 179 B: 68
		4 =>	x"00004CFF", -- R: 255 G: 76 B: 0
		5 =>	x"0041AFFF", -- R: 255 G: 175 B: 65
		6 =>	x"0040AEFF", -- R: 255 G: 174 B: 64
		7 =>	x"000758FF", -- R: 255 G: 88 B: 7
		8 =>	x"000F57FF", -- R: 255 G: 87 B: 15
		9 =>	x"0018B77B", -- R: 123 G: 183 B: 24
		10 =>	x"00000100", -- R: 0 G: 1 B: 0
		11 =>	x"0020B57B", -- R: 123 G: 181 B: 32
		12 =>	x"0000F001", -- R: 1 G: 240 B: 0
		13 =>	x"00000068", -- R: 104 G: 0 B: 0
		14 =>	x"00006500", -- R: 0 G: 101 B: 0
		15 =>	x"0028B37B", -- R: 123 G: 179 B: 40
		16 =>	x"0000B0B3", -- R: 179 G: 176 B: 0
		17 =>	x"007B0070", -- R: 112 G: 0 B: 123
		18 =>	x"008B7700", -- R: 0 G: 119 B: 139
		19 =>	x"00A88B77", -- R: 119 G: 139 B: 168
		20 =>	x"000070B4", -- R: 180 G: 112 B: 0
		21 =>	x"007B0028", -- R: 40 G: 0 B: 123
		22 =>	x"00B47B00", -- R: 0 G: 123 B: 180
		23 =>	x"0000006F", -- R: 111 G: 0 B: 0
		24 =>	x"00BDFC4D", -- R: 77 G: 252 B: 189
		25 =>	x"00A18000", -- R: 0 G: 128 B: 161
		26 =>	x"000C3F0E", -- R: 14 G: 63 B: 12
		27 =>	x"00000009", -- R: 9 G: 0 B: 0
		28 =>	x"00040000", -- R: 0 G: 0 B: 4
		29 =>	x"00518000", -- R: 0 G: 128 B: 81
		30 =>	x"000010B8", -- R: 184 G: 16 B: 0
		31 =>	x"007B0008", -- R: 8 G: 0 B: 123
		32 =>	x"00957700", -- R: 0 G: 119 B: 149
		33 =>	x"00001A00", -- R: 0 G: 26 B: 0
		34 =>	x"00001AB5", -- R: 181 G: 26 B: 0
		35 =>	x"00800000", -- R: 0 G: 0 B: 128
		36 =>	x"0010B87B", -- R: 123 G: 184 B: 16
		37 =>	x"00000895", -- R: 149 G: 8 B: 0
		38 =>	x"00770000", -- R: 0 G: 0 B: 119
		39 =>	x"00DDDDDD", -- R: 221 G: 221 B: 221
		40 =>	x"0000003F", -- R: 63 G: 0 B: 0
		41 =>	x"00E88000", -- R: 0 G: 128 B: 232
		42 =>	x"007B0068", -- R: 104 G: 0 B: 123
		43 =>	x"00AF7B00", -- R: 0 G: 123 B: 175
		44 =>	x"00FDFDFD", -- R: 253 G: 253 B: 253
		45 =>	x"00FDDDDD", -- R: 221 G: 221 B: 253
		46 =>	x"00DDDD30", -- R: 48 G: 221 B: 221
		47 =>	x"00BDFD13", -- R: 19 G: 253 B: 189
		48 =>	x"00F68000", -- R: 0 G: 128 B: 246
		49 =>	x"00DDDD3F", -- R: 63 G: 221 B: 221
		50 =>	x"0040ADFF", -- R: 255 G: 173 B: 64
		51 =>	x"003EABFF", -- R: 255 G: 171 B: 62
		52 =>	x"000E67FF", -- R: 255 G: 103 B: 14
		53 =>	x"00004BFF", -- R: 255 G: 75 B: 0
		54 =>	x"000D56FF", -- R: 255 G: 86 B: 13
		55 =>	x"000556FF", -- R: 255 G: 86 B: 5
		56 =>	x"0038A2FF", -- R: 255 G: 162 B: 56
		57 =>	x"00176DFF", -- R: 255 G: 109 B: 23
		58 =>	x"000F55FF", -- R: 255 G: 85 B: 15
		59 =>	x"001A72FF", -- R: 255 G: 114 B: 26
		60 =>	x"0037A1FF", -- R: 255 G: 161 B: 55
		61 =>	x"003FADFF", -- R: 255 G: 173 B: 63
		62 =>	x"0039A4FF", -- R: 255 G: 164 B: 57
		63 =>	x"000451FF", -- R: 255 G: 81 B: 4
		64 =>	x"003DAAFF", -- R: 255 G: 170 B: 61
		65 =>	x"000D66FF", -- R: 255 G: 102 B: 13
		66 =>	x"000351FF", -- R: 255 G: 81 B: 3
		67 =>	x"001E7BFF", -- R: 255 G: 123 B: 30
		68 =>	x"001877FF", -- R: 255 G: 119 B: 24
		69 =>	x"000F69FF", -- R: 255 G: 105 B: 15
		70 =>	x"00065AFF", -- R: 255 G: 90 B: 6
		71 =>	x"00F2F6FF", -- R: 255 G: 246 B: 242
		72 =>	x"001C77FF", -- R: 255 G: 119 B: 28
		73 =>	x"00F3F7FF", -- R: 255 G: 247 B: 243
		74 =>	x"001A74FF", -- R: 255 G: 116 B: 26
		75 =>	x"00034FFF", -- R: 255 G: 79 B: 3
		76 =>	x"00F6F9FF", -- R: 255 G: 249 B: 246
		77 =>	x"003CA9FF", -- R: 255 G: 169 B: 60
		78 =>	x"003FACFF", -- R: 255 G: 172 B: 63
		79 =>	x"0078A1FF", -- R: 255 G: 161 B: 120
		80 =>	x"00207EFF", -- R: 255 G: 126 B: 32
		81 =>	x"0044B4FF", -- R: 255 G: 180 B: 68
		82 =>	x"002382FF", -- R: 255 G: 130 B: 35
		83 =>	x"006D99FF", -- R: 255 G: 153 B: 109
		84 =>	x"003D0000", -- R: 0 G: 0 B: 61
		85 =>	x"003DEA80", -- R: 128 G: 234 B: 61
		86 =>	x"00000010", -- R: 16 G: 0 B: 0
		87 =>	x"00B87B00", -- R: 0 G: 123 B: 184
		88 =>	x"0068AF7B", -- R: 123 G: 175 B: 104
		89 =>	x"000000D5", -- R: 213 G: 0 B: 0
		90 =>	x"0040F1FF", -- R: 255 G: 241 B: 64
		91 =>	x"000000D4", -- R: 212 G: 0 B: 0
		92 =>	x"000808D6", -- R: 214 G: 8 B: 8
		93 =>	x"000052FF", -- R: 255 G: 82 B: 0
		94 =>	x"00004AFD", -- R: 253 G: 74 B: 0
		95 =>	x"00000CDB", -- R: 219 G: 12 B: 0
		96 =>	x"000A5CFF", -- R: 255 G: 92 B: 10
		97 =>	x"00000DDC", -- R: 220 G: 13 B: 0
		98 =>	x"003CA8FF", -- R: 255 G: 168 B: 60
		99 =>	x"00085AFF", -- R: 255 G: 90 B: 8
		100 =>	x"000B0BD7", -- R: 215 G: 11 B: 11
		101 =>	x"000000D3", -- R: 211 G: 0 B: 0
		102 =>	x"000007D9", -- R: 217 G: 7 B: 0
		103 =>	x"000044FA", -- R: 250 G: 68 B: 0
		104 =>	x"0040EEFF", -- R: 255 G: 238 B: 64
		105 =>	x"0040F5FF", -- R: 255 G: 245 B: 64
		106 =>	x"0040F2FF", -- R: 255 G: 242 B: 64
		107 =>	x"000F0FD7", -- R: 215 G: 15 B: 15
		108 =>	x"000049FF", -- R: 255 G: 73 B: 0
		109 =>	x"000047FC", -- R: 252 G: 71 B: 0
		110 =>	x"0040C9FF", -- R: 255 G: 201 B: 64
		111 =>	x"003BA7FF", -- R: 255 G: 167 B: 59
		112 =>	x"0040ECFF", -- R: 255 G: 236 B: 64
		113 =>	x"00000FDD", -- R: 221 G: 15 B: 0
		114 =>	x"000012DF", -- R: 223 G: 18 B: 0
		115 =>	x"000014E0", -- R: 224 G: 20 B: 0
		116 =>	x"00146CFF", -- R: 255 G: 108 B: 20
		117 =>	x"000041F9", -- R: 249 G: 65 B: 0
		118 =>	x"00004EFF", -- R: 255 G: 78 B: 0
		119 =>	x"000404D6", -- R: 214 G: 4 B: 4
		120 =>	x"0000DEFF", -- R: 255 G: 222 B: 0
		121 =>	x"000010DE", -- R: 222 G: 16 B: 0
		122 =>	x"00004BFE", -- R: 254 G: 75 B: 0
		123 =>	x"0000DFFF", -- R: 255 G: 223 B: 0
		124 =>	x"00004AFF", -- R: 255 G: 74 B: 0
		125 =>	x"0008E2FF", -- R: 255 G: 226 B: 8
		126 =>	x"0040CEFF", -- R: 255 G: 206 B: 64
		127 =>	x"000C60FF", -- R: 255 G: 96 B: 12
		128 =>	x"0000E0FF", -- R: 255 G: 224 B: 0
		129 =>	x"0044B5FF", -- R: 255 G: 181 B: 68
		130 =>	x"000050FF", -- R: 255 G: 80 B: 0
		131 =>	x"000101D5", -- R: 213 G: 1 B: 1
		132 =>	x"000250FF", -- R: 255 G: 80 B: 2
		133 =>	x"0040CDFF", -- R: 255 G: 205 B: 64
		134 =>	x"0041F5FF", -- R: 255 G: 245 B: 65
		135 =>	x"0039F3FF", -- R: 255 G: 243 B: 57
		136 =>	x"000C66FF", -- R: 255 G: 102 B: 12
		137 =>	x"000E6AFF", -- R: 255 G: 106 B: 14
		138 =>	x"0045F7FF", -- R: 255 G: 247 B: 69
		139 =>	x"0045BCFF", -- R: 255 G: 188 B: 69
		140 =>	x"000053FF", -- R: 255 G: 83 B: 0
		141 =>	x"00BDBDF4", -- R: 244 G: 189 B: 189
		142 =>	x"0040C6FF", -- R: 255 G: 198 B: 64
		143 =>	x"000046FF", -- R: 255 G: 70 B: 0
		144 =>	x"005B5BE4", -- R: 228 G: 91 B: 91
		145 =>	x"00002FEF", -- R: 239 G: 47 B: 0
		146 =>	x"000000D2", -- R: 210 G: 0 B: 0
		147 =>	x"000051FF", -- R: 255 G: 81 B: 0
		148 =>	x"002686FF", -- R: 255 G: 134 B: 38
		149 =>	x"000076FF", -- R: 255 G: 118 B: 0
		150 =>	x"0000CDFF", -- R: 255 G: 205 B: 0
		151 =>	x"000087FF", -- R: 255 G: 135 B: 0
		152 =>	x"0004DDFF", -- R: 255 G: 221 B: 4
		153 =>	x"000031F0", -- R: 240 G: 49 B: 0
		154 =>	x"005555E3", -- R: 227 G: 85 B: 85
		155 =>	x"0006DDFF", -- R: 255 G: 221 B: 6
		156 =>	x"0002DEFF", -- R: 255 G: 222 B: 2
		157 =>	x"0004DEFF", -- R: 255 G: 222 B: 4
		158 =>	x"00004CFE", -- R: 254 G: 76 B: 0
		159 =>	x"0000DDFF", -- R: 255 G: 221 B: 0
		160 =>	x"0006DAFF", -- R: 255 G: 218 B: 6
		161 =>	x"0002DDFF", -- R: 255 G: 221 B: 2
		162 =>	x"000040F8", -- R: 248 G: 64 B: 0
		163 =>	x"0040CFFF", -- R: 255 G: 207 B: 64
		164 =>	x"002ED4FF", -- R: 255 G: 212 B: 46
		165 =>	x"0008DDFF", -- R: 255 G: 221 B: 8
		166 =>	x"0028D5FF", -- R: 255 G: 213 B: 40
		167 =>	x"0000D1FF", -- R: 255 G: 209 B: 0
		168 =>	x"0000CCFF", -- R: 255 G: 204 B: 0
		169 =>	x"000083FE", -- R: 254 G: 131 B: 0
		170 =>	x"0012DBFF", -- R: 255 G: 219 B: 18
		171 =>	x"000E69FF", -- R: 255 G: 105 B: 14
		172 =>	x"0025DBFF", -- R: 255 G: 219 B: 37
		173 =>	x"0016DEFF", -- R: 255 G: 222 B: 22
		174 =>	x"000092FF", -- R: 255 G: 146 B: 0
		175 =>	x"001BDCFF", -- R: 255 G: 220 B: 27
		176 =>	x"0018D9FF", -- R: 255 G: 217 B: 24
		177 =>	x"000000D0", -- R: 208 G: 0 B: 0
		178 =>	x"0041BFFF", -- R: 255 G: 191 B: 65
		179 =>	x"003DC6FF", -- R: 255 G: 198 B: 61
		180 =>	x"0040CBFF", -- R: 255 G: 203 B: 64
		181 =>	x"0041CFFF", -- R: 255 G: 207 B: 65
		182 =>	x"0043D6FF", -- R: 255 G: 214 B: 67
		183 =>	x"000044FF", -- R: 255 G: 68 B: 0
		184 =>	x"001E85FF", -- R: 255 G: 133 B: 30
		185 =>	x"00269AFF", -- R: 255 G: 154 B: 38
		186 =>	x"001E8AFF", -- R: 255 G: 138 B: 30
		187 =>	x"000033F1", -- R: 241 G: 51 B: 0
		188 =>	x"004F4FE2", -- R: 226 G: 79 B: 79
		189 =>	x"0040B2FF", -- R: 255 G: 178 B: 64
		190 =>	x"0040AFFF", -- R: 255 G: 175 B: 64
		191 =>	x"0040B1FF", -- R: 255 G: 177 B: 64
		192 =>	x"00C3C3F5", -- R: 245 G: 195 B: 195
		193 =>	x"001871FF", -- R: 255 G: 113 B: 24
		194 =>	x"002688FF", -- R: 255 G: 136 B: 38
		195 =>	x"000202D5", -- R: 213 G: 2 B: 2
		196 =>	x"00F0F0FD", -- R: 253 G: 240 B: 240
		197 =>	x"00CECEF7", -- R: 247 G: 206 B: 206
		198 =>	x"003AA5FF", -- R: 255 G: 165 B: 58
		199 =>	x"0040ACFF", -- R: 255 G: 172 B: 64
		200 =>	x"0040B4FF", -- R: 255 G: 180 B: 64
		201 =>	x"0040B0FF", -- R: 255 G: 176 B: 64
		202 =>	x"0042B2FF", -- R: 255 G: 178 B: 66
		203 =>	x"0042B1FF", -- R: 255 G: 177 B: 66
		204 =>	x"001253F4", -- R: 244 G: 83 B: 18
		205 =>	x"00389EFD", -- R: 253 G: 158 B: 56
		206 =>	x"001268FF", -- R: 255 G: 104 B: 18
		207 =>	x"00002DEE", -- R: 238 G: 45 B: 0
		208 =>	x"003CA7FF", -- R: 255 G: 167 B: 60
		209 =>	x"00006AFF", -- R: 255 G: 106 B: 0
		210 =>	x"00006CFF", -- R: 255 G: 108 B: 0
		211 =>	x"00006BFF", -- R: 255 G: 107 B: 0
		212 =>	x"00FAFAFE", -- R: 254 G: 250 B: 250
		213 =>	x"000069FF", -- R: 255 G: 105 B: 0
		214 =>	x"00005FFF", -- R: 255 G: 95 B: 0
		215 =>	x"00001EE1", -- R: 225 G: 30 B: 0
		216 =>	x"000068FF", -- R: 255 G: 104 B: 0
		217 =>	x"000061FF", -- R: 255 G: 97 B: 0
		218 =>	x"000062FB", -- R: 251 G: 98 B: 0
		219 =>	x"000059FF", -- R: 255 G: 89 B: 0
		220 =>	x"000069FE", -- R: 254 G: 105 B: 0
		221 =>	x"000033E9", -- R: 233 G: 51 B: 0
		222 =>	x"00FDFDFF", -- R: 255 G: 253 B: 253
		223 =>	x"000048FD", -- R: 253 G: 72 B: 0
		224 =>	x"000063FF", -- R: 255 G: 99 B: 0
		225 =>	x"00000FDC", -- R: 220 G: 15 B: 0
		226 =>	x"000059FD", -- R: 253 G: 89 B: 0
		227 =>	x"00D3D3F8", -- R: 248 G: 211 B: 211
		228 =>	x"000055FF", -- R: 255 G: 85 B: 0
		229 =>	x"000051FD", -- R: 253 G: 81 B: 0
		230 =>	x"00006DFF", -- R: 255 G: 109 B: 0
		231 =>	x"000043F0", -- R: 240 G: 67 B: 0
		232 =>	x"00B7B7F3", -- R: 243 G: 183 B: 183
		233 =>	x"00006EFF", -- R: 255 G: 110 B: 0
		234 =>	x"00006BFE", -- R: 254 G: 107 B: 0
		235 =>	x"006060E5", -- R: 229 G: 96 B: 96
		236 =>	x"006464E5", -- R: 229 G: 100 B: 100
		237 =>	x"00000ADA", -- R: 218 G: 10 B: 0
		238 =>	x"007171E8", -- R: 232 G: 113 B: 113
		239 =>	x"00003EEF", -- R: 239 G: 62 B: 0
		240 =>	x"00003BEC", -- R: 236 G: 59 B: 0
		241 =>	x"000039EC", -- R: 236 G: 57 B: 0
		242 =>	x"000030EC", -- R: 236 G: 48 B: 0
		243 =>	x"000011DB", -- R: 219 G: 17 B: 0
		244 =>	x"000034E9", -- R: 233 G: 52 B: 0
		245 =>	x"00002CED", -- R: 237 G: 44 B: 0
		246 =>	x"006666E6", -- R: 230 G: 102 B: 102
		247 =>	x"00008B1F", -- R: 31 G: 139 B: 0
		248 =>	x"00010101", -- R: 1 G: 1 B: 1
		249 =>	x"00B9B9B9", -- R: 185 G: 185 B: 185
		250 =>	x"006C7DF9", -- R: 249 G: 125 B: 108
		251 =>	x"00FFB463", -- R: 99 G: 180 B: 255
		252 =>	x"00001851", -- R: 81 G: 24 B: 0
		253 =>	x"00014D95", -- R: 149 G: 77 B: 1
		254 =>	x"00241CED", -- R: 237 G: 28 B: 36
		others => x"00000000"
	);




begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;