
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);

-- GENERATED BY BC_MEM_PACKER
-- DATE: Mon Jun 06 17:39:44 2016

	signal mem : ram_t := (

--			***** COLOR PALLETE *****


		0 =>	x"00000000", -- R: 0 G: 0 B: 0
		1 =>	x"00008B1F", -- R: 31 G: 139 B: 0
		2 =>	x"00FFFFFF", -- R: 255 G: 255 B: 255
		3 =>	x"00010101", -- R: 1 G: 1 B: 1
		4 =>	x"006C7DF9", -- R: 249 G: 125 B: 108
		5 =>	x"00FFB463", -- R: 99 G: 180 B: 255
		6 =>	x"00B9B9B9", -- R: 185 G: 185 B: 185
		7 =>	x"00001851", -- R: 81 G: 24 B: 0
		8 =>	x"00014D95", -- R: 149 G: 77 B: 1
		9 =>	x"00000000", -- Unused
		10 =>	x"00000000", -- Unused
		11 =>	x"00000000", -- Unused
		12 =>	x"00000000", -- Unused
		13 =>	x"00000000", -- Unused
		14 =>	x"00000000", -- Unused
		15 =>	x"00000000", -- Unused
		16 =>	x"00000000", -- Unused
		17 =>	x"00000000", -- Unused
		18 =>	x"00000000", -- Unused
		19 =>	x"00000000", -- Unused
		20 =>	x"00000000", -- Unused
		21 =>	x"00000000", -- Unused
		22 =>	x"00000000", -- Unused
		23 =>	x"00000000", -- Unused
		24 =>	x"00000000", -- Unused
		25 =>	x"00000000", -- Unused
		26 =>	x"00000000", -- Unused
		27 =>	x"00000000", -- Unused
		28 =>	x"00000000", -- Unused
		29 =>	x"00000000", -- Unused
		30 =>	x"00000000", -- Unused
		31 =>	x"00000000", -- Unused
		32 =>	x"00000000", -- Unused
		33 =>	x"00000000", -- Unused
		34 =>	x"00000000", -- Unused
		35 =>	x"00000000", -- Unused
		36 =>	x"00000000", -- Unused
		37 =>	x"00000000", -- Unused
		38 =>	x"00000000", -- Unused
		39 =>	x"00000000", -- Unused
		40 =>	x"00000000", -- Unused
		41 =>	x"00000000", -- Unused
		42 =>	x"00000000", -- Unused
		43 =>	x"00000000", -- Unused
		44 =>	x"00000000", -- Unused
		45 =>	x"00000000", -- Unused
		46 =>	x"00000000", -- Unused
		47 =>	x"00000000", -- Unused
		48 =>	x"00000000", -- Unused
		49 =>	x"00000000", -- Unused
		50 =>	x"00000000", -- Unused
		51 =>	x"00000000", -- Unused
		52 =>	x"00000000", -- Unused
		53 =>	x"00000000", -- Unused
		54 =>	x"00000000", -- Unused
		55 =>	x"00000000", -- Unused
		56 =>	x"00000000", -- Unused
		57 =>	x"00000000", -- Unused
		58 =>	x"00000000", -- Unused
		59 =>	x"00000000", -- Unused
		60 =>	x"00000000", -- Unused
		61 =>	x"00000000", -- Unused
		62 =>	x"00000000", -- Unused
		63 =>	x"00000000", -- Unused
		64 =>	x"00000000", -- Unused
		65 =>	x"00000000", -- Unused
		66 =>	x"00000000", -- Unused
		67 =>	x"00000000", -- Unused
		68 =>	x"00000000", -- Unused
		69 =>	x"00000000", -- Unused
		70 =>	x"00000000", -- Unused
		71 =>	x"00000000", -- Unused
		72 =>	x"00000000", -- Unused
		73 =>	x"00000000", -- Unused
		74 =>	x"00000000", -- Unused
		75 =>	x"00000000", -- Unused
		76 =>	x"00000000", -- Unused
		77 =>	x"00000000", -- Unused
		78 =>	x"00000000", -- Unused
		79 =>	x"00000000", -- Unused
		80 =>	x"00000000", -- Unused
		81 =>	x"00000000", -- Unused
		82 =>	x"00000000", -- Unused
		83 =>	x"00000000", -- Unused
		84 =>	x"00000000", -- Unused
		85 =>	x"00000000", -- Unused
		86 =>	x"00000000", -- Unused
		87 =>	x"00000000", -- Unused
		88 =>	x"00000000", -- Unused
		89 =>	x"00000000", -- Unused
		90 =>	x"00000000", -- Unused
		91 =>	x"00000000", -- Unused
		92 =>	x"00000000", -- Unused
		93 =>	x"00000000", -- Unused
		94 =>	x"00000000", -- Unused
		95 =>	x"00000000", -- Unused
		96 =>	x"00000000", -- Unused
		97 =>	x"00000000", -- Unused
		98 =>	x"00000000", -- Unused
		99 =>	x"00000000", -- Unused
		100 =>	x"00000000", -- Unused
		101 =>	x"00000000", -- Unused
		102 =>	x"00000000", -- Unused
		103 =>	x"00000000", -- Unused
		104 =>	x"00000000", -- Unused
		105 =>	x"00000000", -- Unused
		106 =>	x"00000000", -- Unused
		107 =>	x"00000000", -- Unused
		108 =>	x"00000000", -- Unused
		109 =>	x"00000000", -- Unused
		110 =>	x"00000000", -- Unused
		111 =>	x"00000000", -- Unused
		112 =>	x"00000000", -- Unused
		113 =>	x"00000000", -- Unused
		114 =>	x"00000000", -- Unused
		115 =>	x"00000000", -- Unused
		116 =>	x"00000000", -- Unused
		117 =>	x"00000000", -- Unused
		118 =>	x"00000000", -- Unused
		119 =>	x"00000000", -- Unused
		120 =>	x"00000000", -- Unused
		121 =>	x"00000000", -- Unused
		122 =>	x"00000000", -- Unused
		123 =>	x"00000000", -- Unused
		124 =>	x"00000000", -- Unused
		125 =>	x"00000000", -- Unused
		126 =>	x"00000000", -- Unused
		127 =>	x"00000000", -- Unused
		128 =>	x"00000000", -- Unused
		129 =>	x"00000000", -- Unused
		130 =>	x"00000000", -- Unused
		131 =>	x"00000000", -- Unused
		132 =>	x"00000000", -- Unused
		133 =>	x"00000000", -- Unused
		134 =>	x"00000000", -- Unused
		135 =>	x"00000000", -- Unused
		136 =>	x"00000000", -- Unused
		137 =>	x"00000000", -- Unused
		138 =>	x"00000000", -- Unused
		139 =>	x"00000000", -- Unused
		140 =>	x"00000000", -- Unused
		141 =>	x"00000000", -- Unused
		142 =>	x"00000000", -- Unused
		143 =>	x"00000000", -- Unused
		144 =>	x"00000000", -- Unused
		145 =>	x"00000000", -- Unused
		146 =>	x"00000000", -- Unused
		147 =>	x"00000000", -- Unused
		148 =>	x"00000000", -- Unused
		149 =>	x"00000000", -- Unused
		150 =>	x"00000000", -- Unused
		151 =>	x"00000000", -- Unused
		152 =>	x"00000000", -- Unused
		153 =>	x"00000000", -- Unused
		154 =>	x"00000000", -- Unused
		155 =>	x"00000000", -- Unused
		156 =>	x"00000000", -- Unused
		157 =>	x"00000000", -- Unused
		158 =>	x"00000000", -- Unused
		159 =>	x"00000000", -- Unused
		160 =>	x"00000000", -- Unused
		161 =>	x"00000000", -- Unused
		162 =>	x"00000000", -- Unused
		163 =>	x"00000000", -- Unused
		164 =>	x"00000000", -- Unused
		165 =>	x"00000000", -- Unused
		166 =>	x"00000000", -- Unused
		167 =>	x"00000000", -- Unused
		168 =>	x"00000000", -- Unused
		169 =>	x"00000000", -- Unused
		170 =>	x"00000000", -- Unused
		171 =>	x"00000000", -- Unused
		172 =>	x"00000000", -- Unused
		173 =>	x"00000000", -- Unused
		174 =>	x"00000000", -- Unused
		175 =>	x"00000000", -- Unused
		176 =>	x"00000000", -- Unused
		177 =>	x"00000000", -- Unused
		178 =>	x"00000000", -- Unused
		179 =>	x"00000000", -- Unused
		180 =>	x"00000000", -- Unused
		181 =>	x"00000000", -- Unused
		182 =>	x"00000000", -- Unused
		183 =>	x"00000000", -- Unused
		184 =>	x"00000000", -- Unused
		185 =>	x"00000000", -- Unused
		186 =>	x"00000000", -- Unused
		187 =>	x"00000000", -- Unused
		188 =>	x"00000000", -- Unused
		189 =>	x"00000000", -- Unused
		190 =>	x"00000000", -- Unused
		191 =>	x"00000000", -- Unused
		192 =>	x"00000000", -- Unused
		193 =>	x"00000000", -- Unused
		194 =>	x"00000000", -- Unused
		195 =>	x"00000000", -- Unused
		196 =>	x"00000000", -- Unused
		197 =>	x"00000000", -- Unused
		198 =>	x"00000000", -- Unused
		199 =>	x"00000000", -- Unused
		200 =>	x"00000000", -- Unused
		201 =>	x"00000000", -- Unused
		202 =>	x"00000000", -- Unused
		203 =>	x"00000000", -- Unused
		204 =>	x"00000000", -- Unused
		205 =>	x"00000000", -- Unused
		206 =>	x"00000000", -- Unused
		207 =>	x"00000000", -- Unused
		208 =>	x"00000000", -- Unused
		209 =>	x"00000000", -- Unused
		210 =>	x"00000000", -- Unused
		211 =>	x"00000000", -- Unused
		212 =>	x"00000000", -- Unused
		213 =>	x"00000000", -- Unused
		214 =>	x"00000000", -- Unused
		215 =>	x"00000000", -- Unused
		216 =>	x"00000000", -- Unused
		217 =>	x"00000000", -- Unused
		218 =>	x"00000000", -- Unused
		219 =>	x"00000000", -- Unused
		220 =>	x"00000000", -- Unused
		221 =>	x"00000000", -- Unused
		222 =>	x"00000000", -- Unused
		223 =>	x"00000000", -- Unused
		224 =>	x"00000000", -- Unused
		225 =>	x"00000000", -- Unused
		226 =>	x"00000000", -- Unused
		227 =>	x"00000000", -- Unused
		228 =>	x"00000000", -- Unused
		229 =>	x"00000000", -- Unused
		230 =>	x"00000000", -- Unused
		231 =>	x"00000000", -- Unused
		232 =>	x"00000000", -- Unused
		233 =>	x"00000000", -- Unused
		234 =>	x"00000000", -- Unused
		235 =>	x"00000000", -- Unused
		236 =>	x"00000000", -- Unused
		237 =>	x"00000000", -- Unused
		238 =>	x"00000000", -- Unused
		239 =>	x"00000000", -- Unused
		240 =>	x"00000000", -- Unused
		241 =>	x"00000000", -- Unused
		242 =>	x"00000000", -- Unused
		243 =>	x"00000000", -- Unused
		244 =>	x"00000000", -- Unused
		245 =>	x"00000000", -- Unused
		246 =>	x"00000000", -- Unused
		247 =>	x"00000000", -- Unused
		248 =>	x"00000000", -- Unused
		249 =>	x"00000000", -- Unused
		250 =>	x"00000000", -- Unused
		251 =>	x"00000000", -- Unused
		252 =>	x"00000000", -- Unused
		253 =>	x"00000000", -- Unused
		254 =>	x"00000000", -- Unused
		
--			***** 8x8 IMAGES *****




--		***** 16x16 IMAGES *****


		255 =>	x"01010101", -- IMG_16x16_bomba
		256 =>	x"01010101",
		257 =>	x"01010101",
		258 =>	x"01010101",
		259 =>	x"01010101",
		260 =>	x"01010101",
		261 =>	x"01020202",
		262 =>	x"01020102",
		263 =>	x"01010101",
		264 =>	x"01030303",
		265 =>	x"02020303",
		266 =>	x"01010101",
		267 =>	x"01010103",
		268 =>	x"03030303",
		269 =>	x"02030303",
		270 =>	x"03010201",
		271 =>	x"01010303",
		272 =>	x"02020303",
		273 =>	x"02030303",
		274 =>	x"03030101",
		275 =>	x"01030302",
		276 =>	x"02030303",
		277 =>	x"03030303",
		278 =>	x"03030301",
		279 =>	x"01030302",
		280 =>	x"02030303",
		281 =>	x"03030303",
		282 =>	x"03030301",
		283 =>	x"03030202",
		284 =>	x"03030303",
		285 =>	x"03030303",
		286 =>	x"03030303",
		287 =>	x"03030202",
		288 =>	x"03030303",
		289 =>	x"03030303",
		290 =>	x"03030303",
		291 =>	x"03030303",
		292 =>	x"03030303",
		293 =>	x"03030303",
		294 =>	x"03030303",
		295 =>	x"03030303",
		296 =>	x"03030303",
		297 =>	x"03030303",
		298 =>	x"03030303",
		299 =>	x"03030303",
		300 =>	x"03030303",
		301 =>	x"03030303",
		302 =>	x"03030303",
		303 =>	x"01030303",
		304 =>	x"03030303",
		305 =>	x"03030303",
		306 =>	x"03030301",
		307 =>	x"01030303",
		308 =>	x"03030303",
		309 =>	x"03030303",
		310 =>	x"03030301",
		311 =>	x"01010303",
		312 =>	x"03030303",
		313 =>	x"03030303",
		314 =>	x"03030101",
		315 =>	x"01010103",
		316 =>	x"03030303",
		317 =>	x"03030303",
		318 =>	x"03010101",
		319 =>	x"01010101", -- IMG_16x16_bomberman
		320 =>	x"01020202",
		321 =>	x"02020201",
		322 =>	x"01010101",
		323 =>	x"01010101",
		324 =>	x"02020202",
		325 =>	x"02020202",
		326 =>	x"01010101",
		327 =>	x"01010101",
		328 =>	x"02040104",
		329 =>	x"04010402",
		330 =>	x"01010101",
		331 =>	x"01010101",
		332 =>	x"02040104",
		333 =>	x"04010402",
		334 =>	x"01010101",
		335 =>	x"01010101",
		336 =>	x"02020202",
		337 =>	x"02020202",
		338 =>	x"01010101",
		339 =>	x"01010101",
		340 =>	x"01020202",
		341 =>	x"02020201",
		342 =>	x"01010101",
		343 =>	x"01010101",
		344 =>	x"01010505",
		345 =>	x"05050101",
		346 =>	x"01010101",
		347 =>	x"01010101",
		348 =>	x"02020505",
		349 =>	x"05050202",
		350 =>	x"01010101",
		351 =>	x"01010102",
		352 =>	x"02050505",
		353 =>	x"05050502",
		354 =>	x"02010101",
		355 =>	x"01010404",
		356 =>	x"02050505",
		357 =>	x"05050502",
		358 =>	x"04040101",
		359 =>	x"01010404",
		360 =>	x"01050505",
		361 =>	x"05050501",
		362 =>	x"04040101",
		363 =>	x"01010101",
		364 =>	x"01050505",
		365 =>	x"05050501",
		366 =>	x"01010101",
		367 =>	x"01010101",
		368 =>	x"01020205",
		369 =>	x"05020201",
		370 =>	x"01010101",
		371 =>	x"01010101",
		372 =>	x"01020201",
		373 =>	x"01020201",
		374 =>	x"01010101",
		375 =>	x"01010101",
		376 =>	x"01040401",
		377 =>	x"01040401",
		378 =>	x"01010101",
		379 =>	x"01010101",
		380 =>	x"01040401",
		381 =>	x"01040401",
		382 =>	x"01010101",
		383 =>	x"02020202", -- IMG_16x16_bombermanBlock
		384 =>	x"02020202",
		385 =>	x"02020202",
		386 =>	x"02020301",
		387 =>	x"06060606",
		388 =>	x"06060606",
		389 =>	x"06060606",
		390 =>	x"06060301",
		391 =>	x"06060606",
		392 =>	x"06060606",
		393 =>	x"06060606",
		394 =>	x"06060301",
		395 =>	x"06060606",
		396 =>	x"06060606",
		397 =>	x"06060606",
		398 =>	x"06060301",
		399 =>	x"06060606",
		400 =>	x"06060606",
		401 =>	x"06060606",
		402 =>	x"06060301",
		403 =>	x"06060606",
		404 =>	x"06060606",
		405 =>	x"06060606",
		406 =>	x"06060301",
		407 =>	x"06060606",
		408 =>	x"06060606",
		409 =>	x"06060606",
		410 =>	x"06060301",
		411 =>	x"06060606",
		412 =>	x"06060606",
		413 =>	x"06060606",
		414 =>	x"06060301",
		415 =>	x"06060606",
		416 =>	x"06060606",
		417 =>	x"06060606",
		418 =>	x"06060301",
		419 =>	x"06060606",
		420 =>	x"06060606",
		421 =>	x"06060606",
		422 =>	x"06060301",
		423 =>	x"06060606",
		424 =>	x"06060606",
		425 =>	x"06060606",
		426 =>	x"06060301",
		427 =>	x"06060606",
		428 =>	x"06060606",
		429 =>	x"06060606",
		430 =>	x"06060301",
		431 =>	x"06060606",
		432 =>	x"06060606",
		433 =>	x"06060606",
		434 =>	x"06060301",
		435 =>	x"06060606",
		436 =>	x"06060606",
		437 =>	x"06060606",
		438 =>	x"06060301",
		439 =>	x"03030303",
		440 =>	x"03030303",
		441 =>	x"03030303",
		442 =>	x"03060301",
		443 =>	x"03030303",
		444 =>	x"03030303",
		445 =>	x"03030303",
		446 =>	x"03030301",
		447 =>	x"03030303", -- IMG_16x16_bombermanBrick
		448 =>	x"03030303",
		449 =>	x"03030303",
		450 =>	x"03030303",
		451 =>	x"03020202",
		452 =>	x"02020202",
		453 =>	x"02020202",
		454 =>	x"02020203",
		455 =>	x"02060606",
		456 =>	x"06060606",
		457 =>	x"06060606",
		458 =>	x"06060603",
		459 =>	x"02060606",
		460 =>	x"06060606",
		461 =>	x"06060606",
		462 =>	x"06060603",
		463 =>	x"02060606",
		464 =>	x"06060606",
		465 =>	x"06060606",
		466 =>	x"06060603",
		467 =>	x"03030303",
		468 =>	x"03030303",
		469 =>	x"03030303",
		470 =>	x"03030303",
		471 =>	x"02020202",
		472 =>	x"02030302",
		473 =>	x"02020202",
		474 =>	x"02020202",
		475 =>	x"06060606",
		476 =>	x"06030206",
		477 =>	x"06060606",
		478 =>	x"06060606",
		479 =>	x"06060606",
		480 =>	x"06030206",
		481 =>	x"06060606",
		482 =>	x"06060606",
		483 =>	x"06060606",
		484 =>	x"06030206",
		485 =>	x"06060606",
		486 =>	x"06060606",
		487 =>	x"03030303",
		488 =>	x"03030303",
		489 =>	x"03030303",
		490 =>	x"03030303",
		491 =>	x"02020202",
		492 =>	x"02020202",
		493 =>	x"02030302",
		494 =>	x"02020202",
		495 =>	x"06060606",
		496 =>	x"06060606",
		497 =>	x"06030206",
		498 =>	x"06060606",
		499 =>	x"06060606",
		500 =>	x"06060606",
		501 =>	x"06030206",
		502 =>	x"06060606",
		503 =>	x"06060606",
		504 =>	x"06060606",
		505 =>	x"06030206",
		506 =>	x"06060606",
		507 =>	x"03030303",
		508 =>	x"03030303",
		509 =>	x"03030303",
		510 =>	x"03030303",
		511 =>	x"03070707", -- IMG_16x16_bombermanDoor
		512 =>	x"07070307",
		513 =>	x"07070707",
		514 =>	x"03030101",
		515 =>	x"07070808",
		516 =>	x"08070307",
		517 =>	x"08080807",
		518 =>	x"07030101",
		519 =>	x"07080807",
		520 =>	x"08070307",
		521 =>	x"08070808",
		522 =>	x"07070101",
		523 =>	x"07080808",
		524 =>	x"08070307",
		525 =>	x"08080808",
		526 =>	x"07070101",
		527 =>	x"07080808",
		528 =>	x"08070307",
		529 =>	x"08080808",
		530 =>	x"07030101",
		531 =>	x"07080803",
		532 =>	x"08070307",
		533 =>	x"08030808",
		534 =>	x"07030101",
		535 =>	x"07080703",
		536 =>	x"07070707",
		537 =>	x"07030708",
		538 =>	x"07030101",
		539 =>	x"07080703",
		540 =>	x"07070707",
		541 =>	x"07030708",
		542 =>	x"07030101",
		543 =>	x"07080803",
		544 =>	x"08070307",
		545 =>	x"08030808",
		546 =>	x"07030101",
		547 =>	x"07080808",
		548 =>	x"08070307",
		549 =>	x"08080808",
		550 =>	x"07030101",
		551 =>	x"07080808",
		552 =>	x"08070307",
		553 =>	x"08080808",
		554 =>	x"07070101",
		555 =>	x"07080807",
		556 =>	x"08070307",
		557 =>	x"08070808",
		558 =>	x"07070101",
		559 =>	x"07070808",
		560 =>	x"08070307",
		561 =>	x"08080807",
		562 =>	x"07030101",
		563 =>	x"03070707",
		564 =>	x"07070307",
		565 =>	x"07070707",
		566 =>	x"03030101",
		567 =>	x"01010101",
		568 =>	x"01010101",
		569 =>	x"01010101",
		570 =>	x"01010101",
		571 =>	x"01010101",
		572 =>	x"01010101",
		573 =>	x"01010101",
		574 =>	x"01010101",
		575 =>	x"01010101", -- IMG_16x16_bombermanEnemie
		576 =>	x"01010101",
		577 =>	x"01010101",
		578 =>	x"01010101",
		579 =>	x"01010101",
		580 =>	x"01010101",
		581 =>	x"01010101",
		582 =>	x"01010101",
		583 =>	x"01010101",
		584 =>	x"03030303",
		585 =>	x"03030303",
		586 =>	x"01010101",
		587 =>	x"01010303",
		588 =>	x"03040404",
		589 =>	x"04040403",
		590 =>	x"03030101",
		591 =>	x"01030304",
		592 =>	x"04040404",
		593 =>	x"04040404",
		594 =>	x"04030301",
		595 =>	x"03030404",
		596 =>	x"04040404",
		597 =>	x"04040404",
		598 =>	x"04040303",
		599 =>	x"03040404",
		600 =>	x"04020204",
		601 =>	x"04020204",
		602 =>	x"04040403",
		603 =>	x"03040404",
		604 =>	x"04030204",
		605 =>	x"04030204",
		606 =>	x"04040403",
		607 =>	x"03040404",
		608 =>	x"04030204",
		609 =>	x"04030204",
		610 =>	x"04040403",
		611 =>	x"03030404",
		612 =>	x"04040404",
		613 =>	x"04040404",
		614 =>	x"04040303",
		615 =>	x"01030404",
		616 =>	x"04040404",
		617 =>	x"04040404",
		618 =>	x"04040301",
		619 =>	x"01030304",
		620 =>	x"04040403",
		621 =>	x"03040404",
		622 =>	x"04030301",
		623 =>	x"01010303",
		624 =>	x"03040404",
		625 =>	x"04040403",
		626 =>	x"03030101",
		627 =>	x"01010101",
		628 =>	x"03030304",
		629 =>	x"04030303",
		630 =>	x"01010101",
		631 =>	x"01010101",
		632 =>	x"01010302",
		633 =>	x"02030101",
		634 =>	x"01010101",
		635 =>	x"01010101",
		636 =>	x"01010303",
		637 =>	x"03030101",
		638 =>	x"01010101",
		639 =>	x"01010101", -- IMG_16x16_pozadinaZeleno
		640 =>	x"01010101",
		641 =>	x"01010101",
		642 =>	x"01010101",
		643 =>	x"01010101",
		644 =>	x"01010101",
		645 =>	x"01010101",
		646 =>	x"01010101",
		647 =>	x"01010101",
		648 =>	x"01010101",
		649 =>	x"01010101",
		650 =>	x"01010101",
		651 =>	x"01010101",
		652 =>	x"01010101",
		653 =>	x"01010101",
		654 =>	x"01010101",
		655 =>	x"01010101",
		656 =>	x"01010101",
		657 =>	x"01010101",
		658 =>	x"01010101",
		659 =>	x"01010101",
		660 =>	x"01010101",
		661 =>	x"01010101",
		662 =>	x"01010101",
		663 =>	x"01010101",
		664 =>	x"01010101",
		665 =>	x"01010101",
		666 =>	x"01010101",
		667 =>	x"01010101",
		668 =>	x"01010101",
		669 =>	x"01010101",
		670 =>	x"01010101",
		671 =>	x"01010101",
		672 =>	x"01010101",
		673 =>	x"01010101",
		674 =>	x"01010101",
		675 =>	x"01010101",
		676 =>	x"01010101",
		677 =>	x"01010101",
		678 =>	x"01010101",
		679 =>	x"01010101",
		680 =>	x"01010101",
		681 =>	x"01010101",
		682 =>	x"01010101",
		683 =>	x"01010101",
		684 =>	x"01010101",
		685 =>	x"01010101",
		686 =>	x"01010101",
		687 =>	x"01010101",
		688 =>	x"01010101",
		689 =>	x"01010101",
		690 =>	x"01010101",
		691 =>	x"01010101",
		692 =>	x"01010101",
		693 =>	x"01010101",
		694 =>	x"01010101",
		695 =>	x"01010101",
		696 =>	x"01010101",
		697 =>	x"01010101",
		698 =>	x"01010101",
		699 =>	x"01010101",
		700 =>	x"01010101",
		701 =>	x"01010101",
		702 =>	x"01010101",



--			***** MAP *****


		703 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		704 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		705 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		706 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		707 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		708 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		709 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		710 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		711 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		712 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		713 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		714 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		715 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		716 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		717 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		718 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		719 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		720 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		721 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		722 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		723 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		724 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		725 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		726 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		727 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		728 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		729 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		730 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		731 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		732 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		733 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		734 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		735 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		736 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		737 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		738 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		739 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		740 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		741 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		742 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		743 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		744 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		745 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		746 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		747 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		748 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		749 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		750 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		751 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		752 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		753 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		754 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		755 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		756 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		757 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		758 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		759 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		760 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		761 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		762 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		763 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		764 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		765 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		766 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		767 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		768 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		769 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		770 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		771 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		772 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		773 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		774 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		775 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		776 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		777 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		778 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		779 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		780 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		781 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		782 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		783 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		784 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		785 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		786 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		787 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		788 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		789 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		790 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		791 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		792 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		793 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		794 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		795 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		796 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		797 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		798 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		799 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		800 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		801 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		802 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		803 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		804 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		805 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		806 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		807 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		808 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		809 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		810 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		811 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		812 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		813 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		814 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		815 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		816 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		817 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		818 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		819 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		820 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		821 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		822 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		823 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		824 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		825 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		826 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		827 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		828 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		829 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		830 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		831 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		832 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		833 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		834 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		835 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		836 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		837 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		838 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		839 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		840 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		841 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		842 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		843 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		844 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		845 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		846 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		847 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		848 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		849 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		850 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		851 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		852 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		853 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		854 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		855 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		856 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		857 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		858 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		859 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		860 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		861 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		862 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		863 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		864 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		865 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		866 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		867 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		868 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		869 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		870 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		871 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		872 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		873 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		874 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		875 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		876 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		877 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		878 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		879 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		880 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		881 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		882 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		883 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		884 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		885 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		886 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		887 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		888 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		889 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		890 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		891 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		892 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		893 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		894 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		895 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		896 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		897 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		898 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		899 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		900 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		901 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		902 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		903 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		904 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		905 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		906 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		907 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		908 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		909 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		910 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		911 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		912 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		913 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		914 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		915 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		916 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		917 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		918 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		919 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		920 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		921 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		922 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		923 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		924 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		925 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		926 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		927 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		928 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		929 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		930 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		931 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		932 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		933 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		934 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		935 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		936 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		937 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		938 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		939 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		940 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		941 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		942 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		943 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		944 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		945 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		946 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		947 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		948 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		949 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		950 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		951 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		952 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		953 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		954 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		955 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		956 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		957 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		958 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		959 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		960 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		961 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		962 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		963 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		964 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		965 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		966 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		967 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		968 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		969 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		970 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		971 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		972 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		973 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		974 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		975 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		976 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		977 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		978 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		979 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		980 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		981 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		982 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		983 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		984 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		985 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		986 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		987 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		988 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		989 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		990 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		991 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		992 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		993 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		994 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		995 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		996 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		997 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		998 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		999 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1000 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1001 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1002 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1003 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1004 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1005 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1006 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1007 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1008 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1009 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1010 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1011 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1012 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1013 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1014 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1015 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1016 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1017 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1018 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1019 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1020 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1021 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1022 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1023 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1024 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1025 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1026 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1027 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1028 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1029 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1030 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1031 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1032 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1033 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1034 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1035 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1036 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1037 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1038 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1039 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1040 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1041 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1042 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1043 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1044 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1045 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1046 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1047 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1048 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1049 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1050 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1051 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1052 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1053 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1054 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1055 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1056 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1057 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1058 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1059 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1060 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1061 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1062 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1063 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1064 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1065 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1066 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1067 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1068 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1069 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1070 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1071 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1072 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1073 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1074 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1075 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1076 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1077 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1078 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1079 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1080 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1081 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1082 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1083 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1084 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1085 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1086 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1087 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1088 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1089 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1090 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1091 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1092 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1093 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1094 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1095 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1096 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1097 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1098 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1099 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1100 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1101 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1102 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1103 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1104 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1105 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1106 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1107 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1108 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1109 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1110 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1111 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1112 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1113 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1114 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1115 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1116 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1117 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1118 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1119 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1120 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1121 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1122 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1123 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1124 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1125 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1126 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1127 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1128 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1129 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1130 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1131 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1132 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1133 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1134 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1135 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1136 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1137 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1138 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1139 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1140 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1141 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1142 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1143 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1144 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1145 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1146 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1147 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1148 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1149 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1150 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1151 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1152 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1153 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1154 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1155 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1156 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1157 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1158 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1159 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1160 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1161 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1162 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1163 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1164 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1165 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1166 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1167 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1168 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1169 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1170 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1171 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1172 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1173 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1174 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1175 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1176 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1177 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1178 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1179 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1180 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1181 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1182 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1183 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1184 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1185 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1186 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1187 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1188 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1189 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1190 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1191 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1192 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1193 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1194 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1195 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1196 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1197 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1198 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1199 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1200 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1201 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1202 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1203 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1204 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1205 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1206 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1207 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1208 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1209 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1210 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1211 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1212 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1213 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1214 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1215 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1216 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1217 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1218 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1219 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1220 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1221 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1222 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1223 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1224 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1225 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1226 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1227 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1228 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1229 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1230 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1231 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1232 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1233 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1234 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1235 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1236 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1237 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1238 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1239 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1240 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1241 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1242 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1243 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1244 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1245 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1246 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1247 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1248 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1249 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1250 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1251 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1252 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1253 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1254 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1255 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1256 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1257 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1258 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1259 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1260 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1261 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1262 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1263 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1264 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1265 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1266 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1267 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1268 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1269 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1270 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1271 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1272 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1273 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1274 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1275 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1276 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1277 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1278 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1279 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1280 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1281 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1282 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1283 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1284 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1285 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1286 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1287 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1288 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1289 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1290 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1291 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1292 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1293 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1294 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1295 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1296 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1297 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1298 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1299 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1300 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1301 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1302 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1303 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1304 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1305 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1306 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1307 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1308 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1309 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1310 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1311 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1312 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1313 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1314 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1315 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1316 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1317 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1318 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1319 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1320 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1321 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1322 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1323 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1324 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1325 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1326 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1327 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1328 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1329 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1330 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1331 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1332 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1333 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1334 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1335 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1336 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1337 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1338 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1339 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1340 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1341 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1342 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1343 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1344 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1345 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1346 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1347 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1348 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1349 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1350 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1351 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1352 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1353 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1354 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1355 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1356 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1357 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1358 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1359 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1360 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1361 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1362 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1363 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1364 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1365 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1366 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1367 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1368 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1369 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1370 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1371 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1372 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1373 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1374 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1375 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1376 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1377 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1378 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1379 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1380 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1381 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1382 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1383 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1384 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1385 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1386 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1387 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1388 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1389 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1390 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1391 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1392 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1393 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1394 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1395 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1396 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1397 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1398 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1399 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1400 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1401 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1402 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1403 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1404 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1405 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1406 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1407 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1408 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1409 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1410 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1411 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1412 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1413 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1414 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1415 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1416 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1417 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1418 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1419 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1420 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1421 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1422 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1423 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1424 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1425 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1426 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1427 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1428 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1429 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1430 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1431 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1432 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1433 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1434 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1435 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1436 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1437 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1438 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1439 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1440 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1441 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1442 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1443 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1444 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1445 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1446 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1447 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1448 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1449 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1450 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1451 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1452 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1453 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1454 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1455 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1456 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1457 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1458 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1459 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1460 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1461 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1462 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1463 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1464 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1465 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1466 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1467 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1468 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1469 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1470 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1471 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1472 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1473 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1474 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1475 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1476 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1477 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1478 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1479 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1480 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1481 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1482 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1483 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1484 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1485 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1486 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1487 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1488 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1489 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1490 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1491 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1492 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1493 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1494 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1495 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1496 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1497 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1498 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1499 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1500 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1501 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1502 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1503 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1504 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1505 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1506 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1507 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1508 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1509 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1510 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1511 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1512 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1513 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1514 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1515 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1516 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1517 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1518 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1519 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1520 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1521 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1522 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1523 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1524 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1525 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1526 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1527 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1528 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1529 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1530 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1531 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1532 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1533 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1534 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1535 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1536 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1537 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1538 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1539 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1540 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1541 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1542 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1543 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1544 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1545 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1546 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1547 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1548 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1549 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1550 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1551 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1552 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1553 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1554 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1555 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1556 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1557 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1558 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1559 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1560 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1561 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1562 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1563 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1564 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1565 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1566 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1567 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1568 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1569 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1570 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1571 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1572 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1573 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1574 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1575 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1576 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1577 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1578 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1579 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1580 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1581 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1582 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1583 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1584 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1585 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1586 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1587 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1588 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1589 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1590 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1591 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1592 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1593 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1594 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1595 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1596 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1597 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1598 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1599 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1600 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1601 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1602 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1603 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1604 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1605 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1606 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1607 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1608 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1609 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1610 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1611 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1612 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1613 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1614 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1615 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1616 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1617 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1618 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1619 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1620 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1621 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1622 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1623 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1624 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1625 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1626 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1627 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1628 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1629 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1630 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1631 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1632 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1633 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1634 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1635 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1636 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1637 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1638 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1639 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1640 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1641 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1642 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1643 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1644 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1645 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1646 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1647 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1648 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1649 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1650 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1651 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1652 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1653 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1654 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1655 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1656 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1657 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1658 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1659 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1660 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1661 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1662 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1663 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1664 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1665 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1666 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1667 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1668 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1669 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1670 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1671 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1672 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1673 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1674 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1675 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1676 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1677 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1678 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1679 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1680 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1681 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1682 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1683 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1684 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1685 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1686 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1687 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1688 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1689 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1690 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1691 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1692 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1693 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1694 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1695 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1696 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1697 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1698 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1699 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1700 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1701 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1702 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1703 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1704 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1705 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1706 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1707 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1708 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1709 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1710 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1711 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1712 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1713 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1714 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1715 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1716 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1717 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1718 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1719 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1720 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1721 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1722 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1723 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1724 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1725 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1726 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1727 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1728 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1729 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1730 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1731 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1732 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1733 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1734 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1735 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1736 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1737 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1738 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1739 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1740 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1741 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1742 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1743 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1744 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1745 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1746 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1747 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1748 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1749 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1750 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1751 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1752 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1753 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1754 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1755 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1756 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1757 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1758 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1759 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1760 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1761 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1762 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1763 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1764 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1765 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1766 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1767 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1768 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1769 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1770 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1771 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1772 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1773 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1774 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1775 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1776 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1777 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1778 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1779 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1780 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1781 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1782 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1783 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1784 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1785 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1786 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1787 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1788 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1789 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1790 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1791 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1792 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1793 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1794 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1795 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1796 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1797 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1798 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1799 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1800 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1801 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1802 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1803 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1804 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1805 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1806 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1807 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1808 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1809 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1810 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1811 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1812 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1813 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1814 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1815 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1816 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1817 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1818 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1819 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1820 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1821 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1822 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1823 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1824 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1825 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1826 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1827 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1828 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1829 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1830 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1831 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1832 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1833 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1834 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1835 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1836 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1837 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1838 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1839 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1840 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1841 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1842 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1843 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1844 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1845 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1846 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1847 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1848 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1849 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1850 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1851 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1852 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1853 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1854 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1855 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1856 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1857 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1858 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1859 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1860 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1861 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1862 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1863 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1864 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1865 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1866 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1867 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1868 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1869 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1870 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1871 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1872 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1873 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1874 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1875 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1876 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1877 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1878 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1879 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1880 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1881 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1882 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1883 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1884 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1885 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1886 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1887 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1888 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1889 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1890 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1891 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1892 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1893 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1894 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1895 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1896 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1897 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1898 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1899 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1900 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1901 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1902 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1903 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1904 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1905 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1906 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1907 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1908 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1909 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1910 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1911 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1912 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1913 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1914 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1915 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1916 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1917 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1918 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1919 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1920 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1921 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1922 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1923 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1924 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1925 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1926 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1927 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1928 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1929 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1930 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1931 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1932 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1933 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1934 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1935 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1936 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1937 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1938 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1939 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1940 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1941 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1942 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1943 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1944 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1945 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1946 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1947 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1948 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1949 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1950 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1951 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1952 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1953 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1954 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1955 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1956 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1957 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1958 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1959 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1960 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1961 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1962 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1963 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1964 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1965 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1966 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1967 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1968 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1969 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1970 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1971 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1972 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1973 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1974 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1975 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1976 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1977 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1978 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1979 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1980 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1981 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1982 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1983 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1984 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1985 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1986 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1987 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1988 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1989 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1990 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1991 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1992 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1993 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1994 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1995 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1996 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1997 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1998 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1999 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2000 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2001 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2002 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2003 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2004 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2005 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2006 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2007 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2008 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2009 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2010 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2011 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2012 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2013 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2014 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2015 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2016 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2017 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2018 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2019 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2020 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2021 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2022 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2023 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2024 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2025 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2026 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2027 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2028 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2029 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2030 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2031 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2032 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2033 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2034 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2035 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2036 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2037 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2038 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2039 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2040 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2041 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2042 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2043 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2044 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2045 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2046 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2047 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2048 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2049 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2050 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2051 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2052 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2053 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2054 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2055 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2056 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2057 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2058 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2059 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2060 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2061 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2062 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2063 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2064 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2065 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2066 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2067 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2068 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2069 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2070 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2071 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2072 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2073 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2074 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2075 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2076 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2077 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2078 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2079 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2080 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2081 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2082 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2083 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2084 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2085 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2086 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2087 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2088 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2089 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2090 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2091 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2092 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2093 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2094 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2095 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2096 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2097 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2098 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2099 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2100 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2101 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2102 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2103 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2104 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2105 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2106 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2107 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2108 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2109 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2110 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2111 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2112 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2113 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2114 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2115 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2116 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2117 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2118 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2119 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2120 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2121 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2122 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2123 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2124 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2125 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2126 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2127 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2128 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2129 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2130 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2131 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2132 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2133 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2134 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2135 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2136 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2137 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2138 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2139 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2140 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2141 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2142 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2143 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2144 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2145 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2146 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2147 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2148 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2149 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2150 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2151 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2152 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2153 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2154 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2155 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2156 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2157 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2158 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2159 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2160 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2161 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2162 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2163 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2164 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2165 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2166 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2167 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2168 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2169 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2170 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2171 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2172 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2173 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2174 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2175 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2176 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2177 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2178 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2179 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2180 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2181 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2182 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2183 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2184 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2185 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2186 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2187 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2188 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2189 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2190 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2191 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2192 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2193 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2194 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2195 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2196 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2197 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2198 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2199 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2200 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2201 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2202 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2203 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2204 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2205 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2206 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2207 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2208 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2209 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2210 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2211 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2212 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2213 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2214 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2215 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2216 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2217 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2218 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2219 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2220 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2221 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2222 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2223 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2224 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2225 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2226 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2227 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2228 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2229 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2230 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2231 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2232 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2233 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2234 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2235 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2236 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2237 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2238 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2239 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2240 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2241 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2242 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2243 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2244 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2245 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2246 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2247 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2248 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2249 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2250 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2251 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2252 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2253 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2254 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2255 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2256 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2257 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2258 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2259 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2260 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2261 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2262 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2263 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2264 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2265 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2266 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2267 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2268 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2269 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2270 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2271 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2272 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2273 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2274 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2275 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2276 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2277 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2278 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2279 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2280 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2281 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2282 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2283 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2284 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2285 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2286 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2287 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2288 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2289 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2290 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2291 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2292 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2293 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2294 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2295 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2296 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2297 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2298 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2299 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2300 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2301 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2302 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2303 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2304 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2305 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2306 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2307 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2308 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2309 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2310 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2311 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2312 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2313 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2314 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2315 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2316 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2317 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2318 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2319 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2320 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2321 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2322 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2323 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2324 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2325 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2326 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2327 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2328 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2329 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2330 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2331 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2332 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2333 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2334 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2335 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2336 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2337 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2338 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2339 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2340 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2341 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2342 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2343 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2344 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2345 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2346 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2347 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2348 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2349 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2350 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2351 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2352 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2353 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2354 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2355 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2356 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2357 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2358 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2359 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2360 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2361 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2362 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2363 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2364 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2365 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2366 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2367 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2368 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2369 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2370 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2371 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2372 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2373 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2374 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2375 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2376 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2377 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2378 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2379 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2380 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2381 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2382 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2383 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2384 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2385 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2386 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2387 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2388 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2389 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2390 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2391 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2392 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2393 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2394 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2395 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2396 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2397 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2398 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2399 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2400 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2401 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2402 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2403 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2404 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2405 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2406 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2407 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2408 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2409 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2410 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2411 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2412 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2413 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2414 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2415 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2416 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2417 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2418 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2419 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2420 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2421 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2422 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2423 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2424 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2425 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2426 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2427 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2428 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2429 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2430 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2431 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2432 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2433 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2434 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2435 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2436 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2437 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2438 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2439 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2440 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2441 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2442 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2443 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2444 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2445 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2446 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2447 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2448 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2449 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2450 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2451 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2452 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2453 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2454 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2455 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2456 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2457 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2458 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2459 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2460 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2461 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2462 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2463 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2464 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2465 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2466 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2467 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2468 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2469 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2470 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2471 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2472 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2473 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2474 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2475 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2476 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2477 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2478 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2479 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2480 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2481 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2482 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2483 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2484 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2485 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2486 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2487 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2488 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2489 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2490 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2491 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2492 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2493 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2494 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2495 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2496 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2497 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2498 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2499 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2500 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2501 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2502 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2503 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2504 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2505 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2506 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2507 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2508 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2509 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2510 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2511 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2512 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2513 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2514 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2515 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2516 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2517 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2518 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2519 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2520 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2521 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2522 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2523 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2524 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2525 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2526 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2527 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2528 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2529 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2530 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2531 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2532 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2533 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2534 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2535 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2536 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2537 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2538 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2539 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2540 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2541 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2542 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2543 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2544 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2545 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2546 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2547 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2548 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2549 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2550 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2551 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2552 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2553 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2554 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2555 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2556 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2557 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2558 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2559 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2560 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2561 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2562 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2563 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2564 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2565 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2566 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2567 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2568 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2569 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2570 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2571 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2572 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2573 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2574 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2575 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2576 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2577 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2578 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2579 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2580 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2581 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2582 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2583 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2584 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2585 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2586 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2587 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2588 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2589 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2590 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2591 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2592 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2593 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2594 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2595 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2596 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2597 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2598 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2599 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2600 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2601 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2602 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2603 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2604 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2605 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2606 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2607 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2608 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2609 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2610 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2611 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2612 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2613 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2614 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2615 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2616 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2617 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2618 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2619 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2620 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2621 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2622 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2623 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2624 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2625 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2626 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2627 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2628 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2629 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2630 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2631 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2632 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2633 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2634 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2635 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2636 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2637 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2638 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2639 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2640 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2641 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2642 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2643 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2644 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2645 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2646 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2647 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2648 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2649 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2650 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2651 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2652 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2653 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2654 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2655 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2656 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2657 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2658 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2659 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2660 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2661 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2662 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2663 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2664 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2665 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2666 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2667 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2668 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2669 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2670 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2671 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2672 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2673 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2674 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2675 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2676 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2677 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2678 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2679 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2680 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2681 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2682 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2683 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2684 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2685 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2686 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2687 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2688 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2689 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2690 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2691 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2692 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2693 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2694 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2695 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2696 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2697 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2698 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2699 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2700 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2701 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2702 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2703 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2704 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2705 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2706 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2707 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2708 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2709 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2710 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2711 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2712 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2713 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2714 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2715 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2716 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2717 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2718 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2719 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2720 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2721 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2722 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2723 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2724 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2725 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2726 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2727 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2728 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2729 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2730 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2731 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2732 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2733 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2734 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2735 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2736 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2737 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2738 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2739 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2740 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2741 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2742 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2743 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2744 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2745 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2746 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2747 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2748 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2749 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2750 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2751 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2752 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2753 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2754 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2755 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2756 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2757 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2758 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2759 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2760 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2761 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2762 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2763 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2764 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2765 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2766 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2767 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2768 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2769 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2770 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2771 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2772 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2773 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2774 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2775 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2776 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2777 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2778 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2779 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2780 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2781 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2782 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2783 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2784 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2785 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2786 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2787 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2788 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2789 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2790 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2791 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2792 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2793 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2794 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2795 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2796 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2797 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2798 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2799 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2800 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2801 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2802 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2803 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2804 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2805 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2806 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2807 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2808 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2809 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2810 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2811 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2812 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2813 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2814 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2815 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2816 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2817 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2818 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2819 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2820 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2821 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2822 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2823 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2824 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2825 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2826 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2827 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2828 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2829 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2830 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2831 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2832 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2833 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2834 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2835 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2836 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2837 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2838 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2839 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2840 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2841 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2842 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2843 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2844 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2845 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2846 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2847 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2848 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2849 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2850 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2851 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2852 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2853 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2854 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2855 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2856 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2857 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2858 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2859 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2860 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2861 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2862 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2863 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2864 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2865 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2866 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2867 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2868 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2869 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2870 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2871 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2872 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2873 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2874 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2875 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2876 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2877 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2878 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2879 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2880 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2881 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2882 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2883 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2884 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2885 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2886 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2887 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2888 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2889 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2890 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2891 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2892 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2893 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2894 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2895 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2896 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2897 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2898 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2899 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2900 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2901 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2902 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2903 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2904 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2905 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2906 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2907 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2908 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2909 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2910 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2911 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2912 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2913 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2914 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2915 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2916 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2917 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2918 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2919 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2920 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2921 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2922 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2923 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2924 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2925 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2926 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2927 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2928 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2929 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2930 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2931 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2932 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2933 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2934 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2935 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2936 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2937 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2938 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2939 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2940 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2941 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2942 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2943 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2944 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2945 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2946 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2947 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2948 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2949 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2950 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2951 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2952 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2953 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2954 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2955 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2956 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2957 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2958 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2959 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2960 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2961 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2962 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2963 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2964 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2965 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2966 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2967 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2968 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2969 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2970 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2971 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2972 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2973 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2974 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2975 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2976 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2977 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2978 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2979 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2980 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2981 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2982 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2983 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2984 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2985 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2986 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2987 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2988 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2989 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2990 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2991 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2992 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2993 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2994 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2995 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2996 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2997 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2998 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2999 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3000 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3001 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3002 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3003 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3004 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3005 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3006 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3007 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3008 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3009 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3010 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3011 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3012 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3013 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3014 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3015 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3016 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3017 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3018 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3019 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3020 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3021 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3022 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3023 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3024 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3025 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3026 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3027 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3028 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3029 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3030 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3031 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3032 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3033 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3034 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3035 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3036 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3037 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3038 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3039 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3040 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3041 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3042 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3043 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3044 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3045 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3046 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3047 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3048 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3049 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3050 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3051 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3052 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3053 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3054 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3055 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3056 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3057 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3058 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3059 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3060 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3061 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3062 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3063 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3064 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3065 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3066 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3067 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3068 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3069 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3070 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3071 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3072 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3073 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3074 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3075 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3076 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3077 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3078 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3079 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3080 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3081 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3082 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3083 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3084 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3085 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3086 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3087 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3088 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3089 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3090 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3091 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3092 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3093 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3094 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3095 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3096 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3097 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3098 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3099 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3100 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3101 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3102 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3103 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3104 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3105 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3106 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3107 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3108 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3109 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3110 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3111 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3112 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3113 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3114 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3115 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3116 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3117 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3118 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3119 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3120 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3121 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3122 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3123 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3124 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3125 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3126 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3127 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3128 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3129 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3130 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3131 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3132 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3133 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3134 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3135 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3136 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3137 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3138 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3139 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3140 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3141 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3142 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3143 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3144 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3145 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3146 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3147 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3148 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3149 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3150 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3151 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3152 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3153 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3154 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3155 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3156 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3157 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3158 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3159 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3160 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3161 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3162 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3163 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3164 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3165 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3166 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3167 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3168 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3169 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3170 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3171 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3172 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3173 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3174 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3175 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3176 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3177 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3178 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3179 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3180 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3181 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3182 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3183 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3184 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3185 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3186 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3187 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3188 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3189 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3190 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3191 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3192 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3193 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3194 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3195 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3196 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3197 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3198 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3199 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3200 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3201 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3202 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3203 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3204 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3205 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3206 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3207 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3208 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3209 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3210 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3211 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3212 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3213 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3214 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3215 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3216 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3217 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3218 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3219 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3220 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3221 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3222 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3223 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3224 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3225 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3226 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3227 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3228 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3229 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3230 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3231 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3232 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3233 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3234 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3235 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3236 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3237 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3238 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3239 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3240 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3241 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3242 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3243 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3244 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3245 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3246 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3247 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3248 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3249 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3250 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3251 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3252 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3253 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3254 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3255 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3256 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3257 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3258 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3259 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3260 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3261 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3262 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3263 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3264 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3265 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3266 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3267 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3268 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3269 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3270 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3271 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3272 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3273 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3274 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3275 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3276 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3277 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3278 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3279 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3280 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3281 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3282 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3283 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3284 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3285 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3286 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3287 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3288 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3289 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3290 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3291 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3292 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3293 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3294 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3295 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3296 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3297 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3298 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3299 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3300 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3301 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3302 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3303 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3304 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3305 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3306 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3307 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3308 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3309 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3310 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3311 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3312 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3313 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3314 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3315 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3316 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3317 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3318 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3319 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3320 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3321 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3322 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3323 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3324 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3325 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3326 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3327 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3328 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3329 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3330 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3331 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3332 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3333 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3334 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3335 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3336 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3337 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3338 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3339 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3340 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3341 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3342 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3343 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3344 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3345 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3346 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3347 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3348 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3349 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3350 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3351 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3352 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3353 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3354 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3355 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3356 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3357 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3358 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3359 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3360 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3361 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3362 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3363 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3364 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3365 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3366 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3367 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3368 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3369 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3370 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3371 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3372 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3373 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3374 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3375 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3376 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3377 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3378 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3379 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3380 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3381 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3382 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3383 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3384 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3385 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3386 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3387 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3388 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3389 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3390 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3391 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3392 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3393 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3394 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3395 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3396 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3397 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3398 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3399 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3400 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3401 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3402 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3403 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3404 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3405 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3406 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3407 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3408 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3409 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3410 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3411 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3412 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3413 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3414 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3415 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3416 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3417 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3418 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3419 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3420 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3421 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3422 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3423 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3424 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3425 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3426 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3427 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3428 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3429 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3430 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3431 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3432 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3433 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3434 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3435 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3436 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3437 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3438 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3439 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3440 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3441 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3442 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3443 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3444 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3445 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3446 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3447 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3448 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3449 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3450 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3451 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3452 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3453 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3454 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3455 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3456 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3457 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3458 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3459 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3460 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3461 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3462 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3463 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3464 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3465 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3466 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3467 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3468 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3469 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3470 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3471 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3472 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3473 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3474 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3475 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3476 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3477 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3478 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3479 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3480 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3481 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3482 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3483 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3484 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3485 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3486 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3487 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3488 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3489 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3490 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3491 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3492 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3493 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3494 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3495 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3496 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3497 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3498 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3499 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3500 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3501 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3502 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3503 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3504 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3505 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3506 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3507 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3508 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3509 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3510 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3511 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3512 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3513 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3514 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3515 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3516 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3517 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3518 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3519 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3520 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3521 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3522 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3523 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3524 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3525 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3526 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3527 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3528 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3529 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3530 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3531 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3532 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3533 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3534 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3535 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3536 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3537 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3538 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3539 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3540 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3541 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3542 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3543 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3544 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3545 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3546 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3547 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3548 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3549 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3550 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3551 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3552 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3553 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3554 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3555 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3556 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3557 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3558 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3559 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3560 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3561 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3562 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3563 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3564 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3565 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3566 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3567 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3568 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3569 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3570 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3571 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3572 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3573 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3574 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3575 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3576 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3577 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3578 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3579 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3580 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3581 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3582 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3583 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3584 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3585 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3586 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3587 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3588 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3589 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3590 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3591 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3592 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3593 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3594 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3595 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3596 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3597 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3598 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3599 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3600 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3601 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3602 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3603 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3604 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3605 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3606 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3607 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3608 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3609 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3610 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3611 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3612 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3613 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3614 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3615 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3616 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3617 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3618 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3619 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3620 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3621 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3622 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3623 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3624 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3625 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3626 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3627 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3628 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3629 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3630 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3631 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3632 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3633 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3634 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3635 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3636 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3637 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3638 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3639 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3640 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3641 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3642 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3643 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3644 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3645 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3646 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3647 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3648 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3649 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3650 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3651 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3652 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3653 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3654 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3655 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3656 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3657 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3658 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3659 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3660 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3661 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3662 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3663 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3664 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3665 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3666 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3667 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3668 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3669 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3670 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3671 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3672 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3673 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3674 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3675 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3676 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3677 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3678 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3679 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3680 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3681 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3682 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3683 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3684 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3685 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3686 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3687 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3688 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3689 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3690 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3691 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3692 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3693 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3694 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3695 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3696 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3697 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3698 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3699 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3700 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3701 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3702 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3703 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3704 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3705 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3706 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3707 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3708 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3709 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3710 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3711 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3712 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3713 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3714 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3715 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3716 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3717 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3718 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3719 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3720 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3721 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3722 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3723 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3724 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3725 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3726 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3727 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3728 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3729 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3730 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3731 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3732 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3733 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3734 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3735 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3736 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3737 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3738 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3739 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3740 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3741 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3742 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3743 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3744 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3745 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3746 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3747 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3748 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3749 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3750 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3751 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3752 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3753 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3754 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3755 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3756 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3757 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3758 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3759 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3760 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3761 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3762 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3763 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3764 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3765 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3766 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3767 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3768 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3769 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3770 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3771 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3772 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3773 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3774 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3775 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3776 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3777 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3778 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3779 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3780 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3781 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3782 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3783 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3784 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3785 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3786 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3787 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3788 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3789 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3790 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3791 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3792 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3793 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3794 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3795 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3796 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3797 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3798 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3799 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3800 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3801 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3802 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3803 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3804 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3805 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3806 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3807 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3808 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3809 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3810 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3811 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3812 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3813 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3814 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3815 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3816 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3817 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3818 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3819 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3820 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3821 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3822 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3823 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3824 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3825 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3826 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3827 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3828 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3829 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3830 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3831 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3832 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3833 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3834 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3835 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3836 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3837 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3838 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3839 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3840 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3841 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3842 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3843 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3844 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3845 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3846 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3847 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3848 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3849 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3850 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3851 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3852 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3853 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3854 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3855 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3856 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3857 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3858 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3859 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3860 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3861 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3862 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3863 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3864 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3865 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3866 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3867 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3868 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3869 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3870 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3871 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3872 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3873 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3874 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3875 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3876 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3877 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3878 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3879 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3880 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3881 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3882 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3883 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3884 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3885 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3886 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3887 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3888 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3889 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3890 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3891 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3892 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3893 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3894 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3895 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3896 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3897 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3898 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3899 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3900 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3901 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3902 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3903 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		3904 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3905 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3906 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3907 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3908 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3909 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3910 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3911 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3912 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3913 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3914 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3915 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3916 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3917 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3918 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3919 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3920 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3921 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3922 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3923 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3924 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3925 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3926 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3927 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3928 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3929 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3930 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3931 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3932 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3933 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3934 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3935 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3936 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3937 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3938 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3939 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3940 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3941 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3942 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3943 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3944 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3945 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3946 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3947 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3948 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3949 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3950 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3951 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3952 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3953 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3954 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3955 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3956 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3957 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3958 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3959 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3960 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3961 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3962 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3963 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3964 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3965 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3966 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3967 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3968 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3969 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3970 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3971 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3972 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3973 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3974 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3975 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3976 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3977 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3978 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3979 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3980 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3981 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3982 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3983 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3984 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3985 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3986 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3987 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3988 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3989 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3990 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3991 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3992 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3993 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3994 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3995 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3996 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3997 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3998 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		3999 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4000 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4001 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4002 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4003 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4004 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4005 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4006 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4007 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4008 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4009 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4010 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4011 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4012 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4013 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4014 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4015 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4016 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4017 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4018 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4019 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4020 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4021 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4022 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4023 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4024 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4025 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4026 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4027 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4028 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4029 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4030 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4031 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4032 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4033 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4034 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4035 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4036 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4037 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4038 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4039 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4040 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4041 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4042 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4043 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4044 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4045 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4046 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4047 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4048 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4049 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4050 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4051 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4052 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4053 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4054 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4055 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4056 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4057 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4058 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4059 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4060 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4061 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4062 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4063 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4064 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4065 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4066 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4067 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4068 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4069 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4070 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4071 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4072 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4073 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4074 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4075 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4076 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4077 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4078 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4079 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4080 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4081 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4082 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4083 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4084 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4085 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4086 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4087 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4088 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4089 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4090 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4091 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4092 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4093 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4094 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4095 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4096 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4097 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4098 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4099 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4100 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4101 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4102 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4103 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4104 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4105 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4106 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4107 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4108 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4109 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4110 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4111 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4112 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4113 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4114 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4115 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4116 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4117 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4118 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4119 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4120 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4121 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4122 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4123 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4124 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4125 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4126 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4127 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4128 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4129 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4130 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4131 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4132 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4133 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4134 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4135 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4136 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4137 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4138 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4139 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4140 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4141 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4142 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4143 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4144 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4145 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4146 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4147 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4148 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4149 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4150 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4151 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4152 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4153 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4154 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4155 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4156 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4157 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4158 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4159 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4160 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4161 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4162 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4163 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4164 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4165 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4166 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4167 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4168 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4169 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4170 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4171 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4172 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4173 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4174 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4175 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4176 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4177 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4178 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4179 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4180 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4181 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4182 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4183 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4184 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4185 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4186 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4187 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4188 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4189 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4190 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4191 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4192 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4193 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4194 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4195 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4196 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4197 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4198 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4199 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4200 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4201 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4202 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4203 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4204 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4205 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4206 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4207 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4208 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4209 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4210 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4211 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4212 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4213 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4214 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4215 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4216 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4217 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4218 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4219 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4220 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4221 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4222 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4223 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4224 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4225 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4226 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4227 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4228 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4229 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4230 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4231 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4232 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4233 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4234 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4235 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4236 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4237 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4238 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4239 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4240 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4241 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4242 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4243 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4244 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4245 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4246 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4247 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4248 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4249 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4250 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4251 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4252 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4253 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4254 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4255 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4256 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4257 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4258 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4259 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4260 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4261 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4262 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4263 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4264 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4265 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4266 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4267 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4268 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4269 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4270 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4271 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4272 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4273 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4274 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4275 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4276 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4277 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4278 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4279 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4280 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4281 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4282 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4283 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4284 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4285 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4286 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4287 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4288 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4289 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4290 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4291 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4292 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4293 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4294 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4295 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4296 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4297 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4298 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4299 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4300 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4301 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4302 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4303 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4304 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4305 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4306 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4307 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4308 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4309 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4310 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4311 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4312 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4313 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4314 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4315 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4316 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4317 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4318 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4319 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4320 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4321 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4322 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4323 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4324 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4325 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4326 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4327 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4328 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4329 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4330 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4331 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4332 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4333 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4334 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4335 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4336 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4337 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4338 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4339 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4340 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4341 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4342 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4343 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4344 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4345 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4346 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4347 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4348 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4349 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4350 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4351 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4352 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4353 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4354 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4355 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4356 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4357 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4358 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4359 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4360 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4361 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4362 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4363 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4364 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4365 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4366 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4367 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4368 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4369 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4370 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4371 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4372 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4373 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4374 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4375 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4376 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4377 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4378 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4379 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4380 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4381 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4382 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4383 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4384 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4385 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4386 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4387 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4388 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4389 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4390 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4391 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4392 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4393 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4394 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4395 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4396 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4397 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4398 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4399 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4400 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4401 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4402 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4403 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4404 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4405 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4406 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4407 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4408 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4409 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4410 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4411 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4412 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4413 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4414 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4415 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4416 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4417 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4418 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4419 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4420 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4421 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4422 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4423 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4424 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4425 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4426 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4427 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4428 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4429 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4430 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4431 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4432 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4433 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4434 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4435 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4436 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4437 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4438 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4439 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4440 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4441 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4442 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4443 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4444 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4445 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4446 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4447 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4448 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4449 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4450 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4451 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4452 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4453 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4454 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4455 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4456 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4457 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4458 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4459 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4460 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4461 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4462 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4463 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4464 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4465 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4466 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4467 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4468 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4469 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4470 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4471 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4472 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4473 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4474 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4475 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4476 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4477 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4478 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4479 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4480 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4481 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4482 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4483 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4484 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4485 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4486 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4487 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4488 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4489 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4490 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4491 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4492 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4493 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4494 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4495 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4496 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4497 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4498 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4499 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4500 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4501 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4502 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4503 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4504 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4505 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4506 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4507 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4508 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4509 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4510 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4511 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4512 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4513 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4514 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4515 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4516 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4517 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4518 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4519 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4520 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4521 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4522 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4523 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4524 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4525 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4526 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4527 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4528 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4529 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4530 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4531 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4532 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4533 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4534 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4535 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4536 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4537 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4538 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4539 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4540 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4541 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4542 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4543 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4544 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4545 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4546 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4547 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4548 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4549 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4550 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4551 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4552 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4553 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4554 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4555 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4556 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4557 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4558 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4559 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4560 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4561 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4562 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4563 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4564 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4565 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4566 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4567 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4568 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4569 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4570 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4571 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4572 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4573 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4574 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4575 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4576 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4577 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4578 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4579 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4580 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4581 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4582 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4583 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4584 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4585 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4586 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4587 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4588 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4589 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4590 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4591 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4592 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4593 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4594 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4595 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4596 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4597 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4598 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4599 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4600 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4601 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4602 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4603 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4604 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4605 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4606 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4607 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4608 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4609 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4610 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4611 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4612 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4613 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4614 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4615 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4616 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4617 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4618 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4619 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4620 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4621 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4622 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4623 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4624 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4625 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4626 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4627 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4628 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4629 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4630 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4631 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4632 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4633 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4634 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4635 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4636 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4637 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4638 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4639 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4640 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4641 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4642 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4643 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4644 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4645 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4646 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4647 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4648 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4649 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4650 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4651 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4652 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4653 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4654 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4655 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4656 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4657 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4658 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4659 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4660 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4661 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4662 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4663 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4664 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4665 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4666 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4667 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4668 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4669 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4670 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4671 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4672 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4673 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4674 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4675 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4676 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4677 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4678 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4679 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4680 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4681 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4682 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4683 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4684 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4685 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4686 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4687 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4688 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4689 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4690 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4691 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4692 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4693 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4694 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4695 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4696 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4697 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4698 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4699 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4700 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4701 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4702 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4703 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4704 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4705 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4706 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4707 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4708 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4709 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4710 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4711 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4712 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4713 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4714 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4715 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4716 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4717 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4718 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4719 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4720 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4721 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4722 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4723 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4724 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4725 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4726 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4727 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4728 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4729 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4730 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4731 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4732 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4733 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4734 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4735 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4736 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4737 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4738 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4739 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4740 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4741 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4742 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4743 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4744 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4745 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4746 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4747 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4748 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4749 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4750 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4751 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4752 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4753 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4754 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4755 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4756 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4757 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4758 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4759 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4760 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4761 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4762 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4763 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4764 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4765 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4766 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4767 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4768 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4769 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4770 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4771 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4772 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4773 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4774 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4775 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4776 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4777 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4778 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4779 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4780 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4781 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4782 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4783 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4784 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4785 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4786 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4787 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4788 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4789 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4790 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4791 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4792 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4793 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4794 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4795 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4796 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4797 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4798 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4799 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4800 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4801 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4802 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4803 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4804 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4805 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4806 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4807 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4808 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4809 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4810 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4811 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4812 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4813 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4814 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4815 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4816 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4817 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4818 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4819 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4820 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4821 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4822 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4823 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4824 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4825 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4826 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4827 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4828 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4829 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4830 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4831 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4832 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4833 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4834 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4835 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4836 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4837 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4838 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4839 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4840 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4841 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4842 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4843 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4844 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4845 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4846 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4847 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4848 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4849 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4850 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4851 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4852 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4853 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4854 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4855 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4856 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4857 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4858 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4859 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4860 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4861 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4862 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4863 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		4864 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4865 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4866 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4867 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4868 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4869 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4870 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4871 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4872 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4873 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4874 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4875 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4876 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4877 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4878 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4879 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4880 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4881 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4882 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4883 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4884 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4885 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4886 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4887 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4888 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4889 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4890 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4891 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4892 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4893 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4894 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4895 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4896 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4897 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4898 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4899 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4900 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4901 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4902 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4903 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4904 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4905 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4906 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4907 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4908 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4909 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4910 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4911 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4912 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4913 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4914 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4915 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4916 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4917 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4918 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4919 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4920 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4921 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4922 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4923 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4924 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4925 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4926 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4927 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4928 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4929 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4930 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4931 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4932 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4933 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4934 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4935 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4936 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4937 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4938 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4939 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4940 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4941 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4942 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4943 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4944 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4945 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4946 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4947 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4948 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4949 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4950 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4951 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4952 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4953 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4954 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4955 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4956 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4957 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4958 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4959 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4960 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4961 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4962 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4963 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4964 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4965 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4966 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4967 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4968 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4969 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4970 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4971 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4972 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4973 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4974 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4975 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4976 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4977 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4978 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4979 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4980 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4981 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4982 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4983 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4984 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4985 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4986 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4987 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4988 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4989 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4990 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4991 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4992 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4993 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4994 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4995 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4996 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4997 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4998 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		4999 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5000 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5001 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5002 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5003 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5004 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5005 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5006 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5007 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5008 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5009 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5010 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5011 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5012 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5013 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5014 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5015 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5016 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5017 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5018 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5019 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5020 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5021 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5022 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5023 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5024 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5025 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5026 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5027 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5028 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5029 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5030 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5031 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5032 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5033 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5034 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5035 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5036 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5037 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5038 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5039 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5040 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5041 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5042 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5043 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5044 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5045 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5046 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5047 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5048 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5049 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5050 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5051 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5052 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5053 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5054 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5055 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5056 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5057 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5058 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5059 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5060 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5061 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5062 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5063 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5064 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5065 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5066 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5067 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5068 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5069 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5070 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5071 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5072 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5073 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5074 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5075 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5076 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5077 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5078 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5079 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5080 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5081 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5082 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5083 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5084 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5085 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5086 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5087 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5088 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5089 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5090 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5091 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5092 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5093 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5094 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5095 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5096 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5097 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5098 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5099 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5100 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5101 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5102 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5103 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5104 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5105 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5106 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5107 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5108 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5109 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5110 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5111 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5112 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5113 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5114 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5115 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5116 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5117 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5118 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5119 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5120 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5121 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5122 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5123 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5124 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5125 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5126 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5127 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5128 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5129 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5130 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5131 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5132 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5133 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5134 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5135 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5136 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5137 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5138 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5139 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5140 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5141 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5142 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5143 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5144 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5145 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5146 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5147 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5148 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5149 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5150 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5151 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5152 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5153 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5154 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5155 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5156 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5157 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5158 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5159 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5160 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5161 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5162 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5163 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5164 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5165 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5166 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5167 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5168 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5169 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5170 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5171 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5172 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5173 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5174 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5175 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5176 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5177 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5178 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5179 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5180 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5181 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5182 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5183 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5184 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5185 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5186 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5187 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5188 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5189 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5190 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5191 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5192 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5193 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5194 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5195 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5196 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5197 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5198 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5199 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5200 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5201 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5202 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5203 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5204 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5205 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5206 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5207 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5208 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5209 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5210 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5211 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5212 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5213 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5214 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5215 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5216 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5217 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5218 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5219 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5220 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5221 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5222 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5223 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5224 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5225 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5226 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5227 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5228 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5229 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5230 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5231 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5232 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5233 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5234 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5235 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5236 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5237 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5238 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5239 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5240 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5241 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5242 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5243 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5244 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5245 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5246 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5247 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5248 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5249 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5250 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5251 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5252 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5253 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5254 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5255 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5256 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5257 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5258 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5259 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5260 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5261 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5262 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5263 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5264 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5265 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5266 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5267 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5268 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5269 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5270 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5271 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5272 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5273 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5274 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5275 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5276 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5277 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5278 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5279 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5280 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5281 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5282 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5283 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5284 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5285 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5286 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5287 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5288 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5289 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5290 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5291 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5292 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5293 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5294 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5295 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5296 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5297 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5298 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5299 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5300 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5301 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5302 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5303 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5304 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5305 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5306 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5307 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5308 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5309 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5310 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5311 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5312 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5313 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5314 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5315 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5316 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5317 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5318 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5319 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5320 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5321 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5322 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5323 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5324 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5325 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5326 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5327 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5328 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5329 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5330 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5331 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5332 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5333 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5334 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5335 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5336 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5337 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5338 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5339 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5340 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5341 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		5342 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5343 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5344 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5345 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5346 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5347 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5348 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5349 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5350 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5351 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5352 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5353 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5354 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5355 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5356 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5357 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5358 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5359 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5360 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5361 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5362 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5363 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5364 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5365 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5366 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5367 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5368 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5369 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5370 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5371 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5372 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5373 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5374 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5375 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5376 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5377 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5378 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5379 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5380 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5381 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5382 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5383 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5384 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5385 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5386 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5387 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5388 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5389 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5390 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5391 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5392 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5393 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5394 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5395 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5396 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5397 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5398 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5399 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5400 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5401 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5402 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5403 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5404 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5405 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5406 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5407 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5408 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5409 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5410 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5411 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5412 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5413 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5414 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5415 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5416 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5417 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5418 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5419 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5420 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5421 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5422 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5423 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5424 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5425 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5426 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5427 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5428 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5429 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5430 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5431 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5432 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5433 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5434 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5435 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5436 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5437 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5438 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5439 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5440 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5441 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5442 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5443 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5444 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5445 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5446 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5447 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5448 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5449 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5450 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5451 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5452 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5453 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5454 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5455 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5456 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5457 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5458 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5459 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5460 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5461 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5462 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5463 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5464 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5465 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5466 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5467 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5468 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5469 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5470 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5471 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5472 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5473 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5474 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5475 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5476 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5477 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5478 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5479 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5480 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5481 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5482 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5483 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5484 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5485 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5486 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5487 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5488 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5489 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5490 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5491 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5492 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5493 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5494 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5495 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5496 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5497 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5498 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5499 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5500 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5501 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		5502 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		others => x"00000000"
	);


begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;