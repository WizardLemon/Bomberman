
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);
-- GENERATED BY BC_MEM_PACKER
-- DATE: Fri May 31 13:35:18 2019

	signal mem : ram_t := (

	
--			***** COLOR PALLETE *****


		0 =>	x"00000000", -- R: 0 G: 0 B: 0
		1 =>	x"00008B1F", -- R: 31 G: 139 B: 0
		2 =>	x"000000D5", -- R: 213 G: 0 B: 0
		3 =>	x"000000D4", -- R: 212 G: 0 B: 0
		4 =>	x"00004DFF", -- R: 255 G: 77 B: 0
		5 =>	x"000041F9", -- R: 249 G: 65 B: 0
		6 =>	x"000052FF", -- R: 255 G: 82 B: 0
		7 =>	x"00004EFF", -- R: 255 G: 78 B: 0
		8 =>	x"000404D6", -- R: 214 G: 4 B: 4
		9 =>	x"0000DEFF", -- R: 255 G: 222 B: 0
		10 =>	x"000010DE", -- R: 222 G: 16 B: 0
		11 =>	x"00004BFF", -- R: 255 G: 75 B: 0
		12 =>	x"00004BFE", -- R: 254 G: 75 B: 0
		13 =>	x"0000DFFF", -- R: 255 G: 223 B: 0
		14 =>	x"00004AFF", -- R: 255 G: 74 B: 0
		15 =>	x"0008E2FF", -- R: 255 G: 226 B: 8
		16 =>	x"0040CEFF", -- R: 255 G: 206 B: 64
		17 =>	x"000C60FF", -- R: 255 G: 96 B: 12
		18 =>	x"0000E0FF", -- R: 255 G: 224 B: 0
		19 =>	x"0044B5FF", -- R: 255 G: 181 B: 68
		20 =>	x"000050FF", -- R: 255 G: 80 B: 0
		21 =>	x"000101D5", -- R: 213 G: 1 B: 1
		22 =>	x"0040F5FF", -- R: 255 G: 245 B: 64
		23 =>	x"0040AEFF", -- R: 255 G: 174 B: 64
		24 =>	x"0041AFFF", -- R: 255 G: 175 B: 65
		25 =>	x"00004CFF", -- R: 255 G: 76 B: 0
		26 =>	x"000808D6", -- R: 214 G: 8 B: 8
		27 =>	x"000250FF", -- R: 255 G: 80 B: 2
		28 =>	x"000049FF", -- R: 255 G: 73 B: 0
		29 =>	x"0040ADFF", -- R: 255 G: 173 B: 64
		30 =>	x"0040CDFF", -- R: 255 G: 205 B: 64
		31 =>	x"0041F5FF", -- R: 255 G: 245 B: 65
		32 =>	x"0039F3FF", -- R: 255 G: 243 B: 57
		33 =>	x"000C66FF", -- R: 255 G: 102 B: 12
		34 =>	x"000E6AFF", -- R: 255 G: 106 B: 14
		35 =>	x"0045F7FF", -- R: 255 G: 247 B: 69
		36 =>	x"0045BCFF", -- R: 255 G: 188 B: 69
		37 =>	x"000012DF", -- R: 223 G: 18 B: 0
		38 =>	x"000053FF", -- R: 255 G: 83 B: 0
		39 =>	x"00BDBDF4", -- R: 244 G: 189 B: 189
		40 =>	x"000014E0", -- R: 224 G: 20 B: 0
		41 =>	x"0040C6FF", -- R: 255 G: 198 B: 64
		42 =>	x"000046FF", -- R: 255 G: 70 B: 0
		43 =>	x"005B5BE4", -- R: 228 G: 91 B: 91
		44 =>	x"00002FEF", -- R: 239 G: 47 B: 0
		45 =>	x"000000D2", -- R: 210 G: 0 B: 0
		46 =>	x"000051FF", -- R: 255 G: 81 B: 0
		47 =>	x"002686FF", -- R: 255 G: 134 B: 38
		48 =>	x"000076FF", -- R: 255 G: 118 B: 0
		49 =>	x"0000CDFF", -- R: 255 G: 205 B: 0
		50 =>	x"000087FF", -- R: 255 G: 135 B: 0
		51 =>	x"0004DDFF", -- R: 255 G: 221 B: 4
		52 =>	x"000031F0", -- R: 240 G: 49 B: 0
		53 =>	x"005555E3", -- R: 227 G: 85 B: 85
		54 =>	x"00020000", -- R: 0 G: 0 B: 2
		55 =>	x"00000F00", -- R: 0 G: 15 B: 0
		56 =>	x"0000000C", -- R: 12 G: 0 B: 0
		57 =>	x"00FDFDFD", -- R: 253 G: 253 B: 253
		58 =>	x"00FD4144", -- R: 68 G: 65 B: 253
		59 =>	x"00564958", -- R: 88 G: 73 B: 86
		60 =>	x"00455F4C", -- R: 76 G: 95 B: 69
		61 =>	x"00414E47", -- R: 71 G: 78 B: 65
		62 =>	x"003D656E", -- R: 110 G: 101 B: 61
		63 =>	x"0000FDFD", -- R: 253 G: 253 B: 0
		64 =>	x"00FDFD00", -- R: 0 G: 253 B: 253
		65 =>	x"0000C551", -- R: 81 G: 197 B: 0
		66 =>	x"001A1A34", -- R: 52 G: 26 B: 26
		67 =>	x"0037000D", -- R: 13 G: 0 B: 55
		68 =>	x"006F6F6C", -- R: 108 G: 111 B: 111
		69 =>	x"00735C41", -- R: 65 G: 92 B: 115
		70 =>	x"00647669", -- R: 105 G: 118 B: 100
		71 =>	x"00736F72", -- R: 114 G: 111 B: 115
		72 =>	x"00203230", -- R: 48 G: 50 B: 32
		73 =>	x"0031375C", -- R: 92 G: 55 B: 49
		74 =>	x"00C7511A", -- R: 26 G: 81 B: 199
		75 =>	x"00183237", -- R: 55 G: 50 B: 24
		76 =>	x"00000D48", -- R: 72 G: 13 B: 0
		77 =>	x"00BC9A00", -- R: 0 G: 154 B: 188
		78 =>	x"00F8BC9A", -- R: 154 G: 188 B: 248
		79 =>	x"00007857", -- R: 87 G: 120 B: 0
		80 =>	x"00355081", -- R: 129 G: 80 B: 53
		81 =>	x"00414456", -- R: 86 G: 68 B: 65
		82 =>	x"0049534F", -- R: 79 G: 83 B: 73
		83 =>	x"00525F32", -- R: 50 G: 95 B: 82
		84 =>	x"00303137", -- R: 55 G: 49 B: 48
		85 =>	x"005F4449", -- R: 73 G: 68 B: 95
		86 =>	x"00523D43", -- R: 67 G: 61 B: 82
		87 =>	x"003A5C50", -- R: 80 G: 92 B: 58
		88 =>	x"00726F67", -- R: 103 G: 111 B: 114
		89 =>	x"0072616D", -- R: 109 G: 97 B: 114
		90 =>	x"00204669", -- R: 105 G: 70 B: 32
		91 =>	x"006C6573", -- R: 115 G: 101 B: 108
		92 =>	x"00202878", -- R: 120 G: 40 B: 32
		93 =>	x"00383629", -- R: 41 G: 54 B: 56
		94 =>	x"005C496E", -- R: 110 G: 73 B: 92
		95 =>	x"0074656C", -- R: 108 G: 101 B: 116
		96 =>	x"00535754", -- R: 84 G: 87 B: 83
		97 =>	x"000000C1", -- R: 193 G: 0 B: 0
		98 =>	x"00511A1E", -- R: 30 G: 26 B: 81
		99 =>	x"00743700", -- R: 0 G: 55 B: 116
		100 =>	x"0009F88D", -- R: 141 G: 248 B: 9
		101 =>	x"009600B8", -- R: 184 G: 0 B: 150
		102 =>	x"00785735", -- R: 53 G: 87 B: 120
		103 =>	x"00508100", -- R: 0 G: 129 B: 80
		104 =>	x"00000002", -- R: 2 G: 0 B: 0
		105 =>	x"00430000", -- R: 0 G: 0 B: 67
		106 =>	x"00000B00", -- R: 0 G: 11 B: 0
		107 =>	x"000000FD", -- R: 253 G: 0 B: 0
		108 =>	x"00001100", -- R: 0 G: 17 B: 0
		109 =>	x"00001179", -- R: 121 G: 17 B: 0
		110 =>	x"00370000", -- R: 0 G: 0 B: 55
		111 =>	x"0018AC9A", -- R: 154 G: 172 B: 24
		112 =>	x"0000C400", -- R: 0 G: 196 B: 0
		113 =>	x"00960000", -- R: 0 G: 0 B: 150
		114 =>	x"00DDDDDD", -- R: 221 G: 221 B: 221
		115 =>	x"00DDDD36", -- R: 54 G: 221 B: 221
		116 =>	x"00000036", -- R: 54 G: 0 B: 0
		117 =>	x"00243700", -- R: 0 G: 55 B: 36
		118 =>	x"000018AC", -- R: 172 G: 24 B: 0
		119 =>	x"009A0070", -- R: 112 G: 0 B: 154
		120 =>	x"00B99A00", -- R: 0 G: 154 B: 185
		121 =>	x"00340000", -- R: 0 G: 0 B: 52
		122 =>	x"00342637", -- R: 55 G: 38 B: 52
		123 =>	x"00000018", -- R: 24 G: 0 B: 0
		124 =>	x"00AC9A00", -- R: 0 G: 154 B: 172
		125 =>	x"0070B99A", -- R: 154 G: 185 B: 112
		126 =>	x"00FDDDDD", -- R: 221 G: 221 B: 253
		127 =>	x"00DDDD87", -- R: 135 G: 221 B: 221
		128 =>	x"00511B59", -- R: 89 G: 27 B: 81
		129 =>	x"003A3700", -- R: 0 G: 55 B: 58
		130 =>	x"00FFFFFF", -- R: 255 G: 255 B: 255
		131 =>	x"0040CFFF", -- R: 255 G: 207 B: 64
		132 =>	x"002ED4FF", -- R: 255 G: 212 B: 46
		133 =>	x"0004DEFF", -- R: 255 G: 222 B: 4
		134 =>	x"0008DDFF", -- R: 255 G: 221 B: 8
		135 =>	x"0028D5FF", -- R: 255 G: 213 B: 40
		136 =>	x"0000D1FF", -- R: 255 G: 209 B: 0
		137 =>	x"0000CCFF", -- R: 255 G: 204 B: 0
		138 =>	x"000083FE", -- R: 254 G: 131 B: 0
		139 =>	x"0002DEFF", -- R: 255 G: 222 B: 2
		140 =>	x"0006DDFF", -- R: 255 G: 221 B: 6
		141 =>	x"0012DBFF", -- R: 255 G: 219 B: 18
		142 =>	x"000E69FF", -- R: 255 G: 105 B: 14
		143 =>	x"0025DBFF", -- R: 255 G: 219 B: 37
		144 =>	x"0016DEFF", -- R: 255 G: 222 B: 22
		145 =>	x"000092FF", -- R: 255 G: 146 B: 0
		146 =>	x"001BDCFF", -- R: 255 G: 220 B: 27
		147 =>	x"0018D9FF", -- R: 255 G: 217 B: 24
		148 =>	x"000000D0", -- R: 208 G: 0 B: 0
		149 =>	x"0041BFFF", -- R: 255 G: 191 B: 65
		150 =>	x"003DC6FF", -- R: 255 G: 198 B: 61
		151 =>	x"0040CBFF", -- R: 255 G: 203 B: 64
		152 =>	x"0041CFFF", -- R: 255 G: 207 B: 65
		153 =>	x"0043D6FF", -- R: 255 G: 214 B: 67
		154 =>	x"000044FF", -- R: 255 G: 68 B: 0
		155 =>	x"001E85FF", -- R: 255 G: 133 B: 30
		156 =>	x"00269AFF", -- R: 255 G: 154 B: 38
		157 =>	x"001E8AFF", -- R: 255 G: 138 B: 30
		158 =>	x"000033F1", -- R: 241 G: 51 B: 0
		159 =>	x"004F4FE2", -- R: 226 G: 79 B: 79
		160 =>	x"003AA5FF", -- R: 255 G: 165 B: 58
		161 =>	x"00004AFD", -- R: 253 G: 74 B: 0
		162 =>	x"0040AFFF", -- R: 255 G: 175 B: 64
		163 =>	x"003BA7FF", -- R: 255 G: 167 B: 59
		164 =>	x"0040ACFF", -- R: 255 G: 172 B: 64
		165 =>	x"0040B1FF", -- R: 255 G: 177 B: 64
		166 =>	x"0040B2FF", -- R: 255 G: 178 B: 64
		167 =>	x"0040B4FF", -- R: 255 G: 180 B: 64
		168 =>	x"0040B0FF", -- R: 255 G: 176 B: 64
		169 =>	x"0042B2FF", -- R: 255 G: 178 B: 66
		170 =>	x"0042B1FF", -- R: 255 G: 177 B: 66
		171 =>	x"003EABFF", -- R: 255 G: 171 B: 62
		172 =>	x"001253F4", -- R: 244 G: 83 B: 18
		173 =>	x"00389EFD", -- R: 253 G: 158 B: 56
		174 =>	x"001268FF", -- R: 255 G: 104 B: 18
		175 =>	x"003CA8FF", -- R: 255 G: 168 B: 60
		176 =>	x"00002DEE", -- R: 238 G: 45 B: 0
		177 =>	x"003CA7FF", -- R: 255 G: 167 B: 60
		178 =>	x"001E7BFF", -- R: 255 G: 123 B: 30
		179 =>	x"000000D3", -- R: 211 G: 0 B: 0
		180 =>	x"00006AFF", -- R: 255 G: 106 B: 0
		181 =>	x"00006CFF", -- R: 255 G: 108 B: 0
		182 =>	x"00006BFF", -- R: 255 G: 107 B: 0
		183 =>	x"00FAFAFE", -- R: 254 G: 250 B: 250
		184 =>	x"000069FF", -- R: 255 G: 105 B: 0
		185 =>	x"00005FFF", -- R: 255 G: 95 B: 0
		186 =>	x"00001EE1", -- R: 225 G: 30 B: 0
		187 =>	x"000068FF", -- R: 255 G: 104 B: 0
		188 =>	x"000061FF", -- R: 255 G: 97 B: 0
		189 =>	x"000062FB", -- R: 251 G: 98 B: 0
		190 =>	x"000059FF", -- R: 255 G: 89 B: 0
		191 =>	x"000069FE", -- R: 254 G: 105 B: 0
		192 =>	x"000033E9", -- R: 233 G: 51 B: 0
		193 =>	x"00000DDC", -- R: 220 G: 13 B: 0
		194 =>	x"00FDFDFF", -- R: 255 G: 253 B: 253
		195 =>	x"000048FD", -- R: 253 G: 72 B: 0
		196 =>	x"000063FF", -- R: 255 G: 99 B: 0
		197 =>	x"00000FDC", -- R: 220 G: 15 B: 0
		198 =>	x"000059FD", -- R: 253 G: 89 B: 0
		199 =>	x"00000CDB", -- R: 219 G: 12 B: 0
		200 =>	x"00D3D3F8", -- R: 248 G: 211 B: 211
		201 =>	x"000055FF", -- R: 255 G: 85 B: 0
		202 =>	x"000047FC", -- R: 252 G: 71 B: 0
		203 =>	x"000051FD", -- R: 253 G: 81 B: 0
		204 =>	x"00006DFF", -- R: 255 G: 109 B: 0
		205 =>	x"000043F0", -- R: 240 G: 67 B: 0
		206 =>	x"00000FDD", -- R: 221 G: 15 B: 0
		207 =>	x"00B7B7F3", -- R: 243 G: 183 B: 183
		208 =>	x"007171E8", -- R: 232 G: 113 B: 113
		209 =>	x"00003EEF", -- R: 239 G: 62 B: 0
		210 =>	x"00003BEC", -- R: 236 G: 59 B: 0
		211 =>	x"000039EC", -- R: 236 G: 57 B: 0
		212 =>	x"000030EC", -- R: 236 G: 48 B: 0
		213 =>	x"000011DB", -- R: 219 G: 17 B: 0
		214 =>	x"000034E9", -- R: 233 G: 52 B: 0
		215 =>	x"00002CED", -- R: 237 G: 44 B: 0
		216 =>	x"006666E6", -- R: 230 G: 102 B: 102
		217 =>	x"00010101", -- R: 1 G: 1 B: 1
		218 =>	x"00B9B9B9", -- R: 185 G: 185 B: 185
		219 =>	x"006C7DF9", -- R: 249 G: 125 B: 108
		220 =>	x"00FFB463", -- R: 99 G: 180 B: 255
		221 =>	x"00001851", -- R: 81 G: 24 B: 0
		222 =>	x"00014D95", -- R: 149 G: 77 B: 1
		223 =>	x"00241CED", -- R: 237 G: 28 B: 36
		224 =>	x"00000000", -- Unused
		225 =>	x"00000000", -- Unused
		226 =>	x"00000000", -- Unused
		227 =>	x"00000000", -- Unused
		228 =>	x"00000000", -- Unused
		229 =>	x"00000000", -- Unused
		230 =>	x"00000000", -- Unused
		231 =>	x"00000000", -- Unused
		232 =>	x"00000000", -- Unused
		233 =>	x"00000000", -- Unused
		234 =>	x"00000000", -- Unused
		235 =>	x"00000000", -- Unused
		236 =>	x"00000000", -- Unused
		237 =>	x"00000000", -- Unused
		238 =>	x"00000000", -- Unused
		239 =>	x"00000000", -- Unused
		240 =>	x"00000000", -- Unused
		241 =>	x"00000000", -- Unused
		242 =>	x"00000000", -- Unused
		243 =>	x"00000000", -- Unused
		244 =>	x"00000000", -- Unused
		245 =>	x"00000000", -- Unused
		246 =>	x"00000000", -- Unused
		247 =>	x"00000000", -- Unused
		248 =>	x"00000000", -- Unused
		249 =>	x"00000000", -- Unused
		250 =>	x"00000000", -- Unused
		251 =>	x"00000000", -- Unused
		252 =>	x"00000000", -- Unused
		253 =>	x"00000000", -- Unused
		254 =>	x"00000000", -- Unused
	
--			***** 16x16 IMAGES *****


		255 =>	x"01010101", -- IMG_16x16_3end_up
		256 =>	x"02020202",
		257 =>	x"02020202",
		258 =>	x"02020101",
		259 =>	x"01010101",
		260 =>	x"03040506",
		261 =>	x"07020404",
		262 =>	x"03020801",
		263 =>	x"01010103",
		264 =>	x"04090909",
		265 =>	x"09090904",
		266 =>	x"04030101",
		267 =>	x"0101010A",
		268 =>	x"0B090909",
		269 =>	x"09090909",
		270 =>	x"040C0801",
		271 =>	x"01010103",
		272 =>	x"0B09090D",
		273 =>	x"09090909",
		274 =>	x"0E030101",
		275 =>	x"0101010A",
		276 =>	x"0B09090D",
		277 =>	x"09090909",
		278 =>	x"0E030801",
		279 =>	x"01010103",
		280 =>	x"0409090F",
		281 =>	x"09090909",
		282 =>	x"100C0801",
		283 =>	x"01010106",
		284 =>	x"11090912",
		285 =>	x"09090909",
		286 =>	x"0E030801",
		287 =>	x"0101010A",
		288 =>	x"0B090909",
		289 =>	x"09090909",
		290 =>	x"0E0C0801",
		291 =>	x"0101010A",
		292 =>	x"04090909",
		293 =>	x"09090909",
		294 =>	x"09040801",
		295 =>	x"0101010A",
		296 =>	x"11090909",
		297 =>	x"09090909",
		298 =>	x"09030101",
		299 =>	x"0101010A",
		300 =>	x"13090909",
		301 =>	x"09090909",
		302 =>	x"09020101",
		303 =>	x"0101010A",
		304 =>	x"0B090909",
		305 =>	x"09090909",
		306 =>	x"04040801",
		307 =>	x"01010102",
		308 =>	x"14090909",
		309 =>	x"09090909",
		310 =>	x"0E0C0801",
		311 =>	x"01010103",
		312 =>	x"0B090909",
		313 =>	x"09090909",
		314 =>	x"0E030801",
		315 =>	x"0101010A",
		316 =>	x"11090909",
		317 =>	x"09090909",
		318 =>	x"04040201",
		319 =>	x"01011502", -- IMG_16x16_3intersection
		320 =>	x"04161616",
		321 =>	x"16161617",
		322 =>	x"07020101",
		323 =>	x"01010204",
		324 =>	x"18161616",
		325 =>	x"16161616",
		326 =>	x"19030101",
		327 =>	x"1A020C04",
		328 =>	x"16161616",
		329 =>	x"16161616",
		330 =>	x"1B04021A",
		331 =>	x"030E040E",
		332 =>	x"16161616",
		333 =>	x"16161616",
		334 =>	x"1C040403",
		335 =>	x"1D1D1E16",
		336 =>	x"16161616",
		337 =>	x"16161616",
		338 =>	x"16161616",
		339 =>	x"16161616",
		340 =>	x"16161616",
		341 =>	x"16161616",
		342 =>	x"16161616",
		343 =>	x"16161616",
		344 =>	x"16161616",
		345 =>	x"16161616",
		346 =>	x"16161616",
		347 =>	x"1F201616",
		348 =>	x"16161616",
		349 =>	x"1616161F",
		350 =>	x"20161F1F",
		351 =>	x"16161616",
		352 =>	x"16161616",
		353 =>	x"16161616",
		354 =>	x"16161616",
		355 =>	x"16161616",
		356 =>	x"16161616",
		357 =>	x"16161616",
		358 =>	x"16161616",
		359 =>	x"16161616",
		360 =>	x"16161616",
		361 =>	x"16161616",
		362 =>	x"16161616",
		363 =>	x"21161616",
		364 =>	x"16161616",
		365 =>	x"16161616",
		366 =>	x"16161721",
		367 =>	x"0604040B",
		368 =>	x"22161623",
		369 =>	x"16161616",
		370 =>	x"24040B06",
		371 =>	x"02252604",
		372 =>	x"04161616",
		373 =>	x"16231616",
		374 =>	x"04042502",
		375 =>	x"01270204",
		376 =>	x"04161616",
		377 =>	x"16161616",
		378 =>	x"04282701",
		379 =>	x"0101020A",
		380 =>	x"04291616",
		381 =>	x"16161616",
		382 =>	x"2A020101",
		383 =>	x"01010101", -- IMG_16x16_3middle_horizontal
		384 =>	x"01010101",
		385 =>	x"01010101",
		386 =>	x"01010101",
		387 =>	x"01010101",
		388 =>	x"01010101",
		389 =>	x"01010101",
		390 =>	x"01010101",
		391 =>	x"2B2B0101",
		392 =>	x"012B2B2B",
		393 =>	x"2B012B2B",
		394 =>	x"0101012B",
		395 =>	x"2C2D022C",
		396 =>	x"2C2C2C2C",
		397 =>	x"2E2D2C2D",
		398 =>	x"2C2D022C",
		399 =>	x"2F2A0E12",
		400 =>	x"12123031",
		401 =>	x"12121212",
		402 =>	x"1212322F",
		403 =>	x"12121212",
		404 =>	x"12121212",
		405 =>	x"12121212",
		406 =>	x"12121233",
		407 =>	x"12121212",
		408 =>	x"12121212",
		409 =>	x"12121212",
		410 =>	x"12121212",
		411 =>	x"12121212",
		412 =>	x"12121212",
		413 =>	x"12121212",
		414 =>	x"12121212",
		415 =>	x"12121212",
		416 =>	x"12121212",
		417 =>	x"12121212",
		418 =>	x"12121212",
		419 =>	x"12121212",
		420 =>	x"12121212",
		421 =>	x"12121212",
		422 =>	x"12121212",
		423 =>	x"12121212",
		424 =>	x"12121212",
		425 =>	x"12121212",
		426 =>	x"12121212",
		427 =>	x"12121212",
		428 =>	x"12121212",
		429 =>	x"12121212",
		430 =>	x"12121212",
		431 =>	x"06121212",
		432 =>	x"12121212",
		433 =>	x"12121212",
		434 =>	x"12041212",
		435 =>	x"2E2D342E",
		436 =>	x"022D2E34",
		437 =>	x"2D342D2D",
		438 =>	x"342D3434",
		439 =>	x"02353535",
		440 =>	x"01013535",
		441 =>	x"35353501",
		442 =>	x"35010101",
		443 =>	x"01010101",
		444 =>	x"01010101",
		445 =>	x"01010101",
		446 =>	x"01010101",
		447 =>	x"36373800", -- IMG_16x16_4end_up
		448 =>	x"393A3B3C",
		449 =>	x"3D3E3F40",
		450 =>	x"00414243",
		451 =>	x"44454647",
		452 =>	x"48493F40",
		453 =>	x"4A4B4C4D",
		454 =>	x"4E4F5000",
		455 =>	x"51525354",
		456 =>	x"55565758",
		457 =>	x"595A5B5C",
		458 =>	x"5D5E5F60",
		459 =>	x"00006162",
		460 =>	x"6364654D",
		461 =>	x"66676800",
		462 =>	x"696A6B39",
		463 =>	x"00000000",
		464 =>	x"00000000",
		465 =>	x"00000000",
		466 =>	x"00000000",
		467 =>	x"00000000",
		468 =>	x"00000000",
		469 =>	x"00000000",
		470 =>	x"00000000",
		471 =>	x"00000000",
		472 =>	x"006C6D6E",
		473 =>	x"6F707100",
		474 =>	x"00000000",
		475 =>	x"00000000",
		476 =>	x"00000000",
		477 =>	x"00000000",
		478 =>	x"00000000",
		479 =>	x"00000000",
		480 =>	x"00000000",
		481 =>	x"00000000",
		482 =>	x"00000000",
		483 =>	x"00000000",
		484 =>	x"00000000",
		485 =>	x"00000000",
		486 =>	x"00000000",
		487 =>	x"00000000",
		488 =>	x"00000000",
		489 =>	x"00000000",
		490 =>	x"00000000",
		491 =>	x"00000000",
		492 =>	x"00000000",
		493 =>	x"00000000",
		494 =>	x"00000000",
		495 =>	x"72727374",
		496 =>	x"75767778",
		497 =>	x"797A7B7C",
		498 =>	x"7D000000",
		499 =>	x"72727272",
		500 =>	x"72727272",
		501 =>	x"72727272",
		502 =>	x"72727272",
		503 =>	x"72727272",
		504 =>	x"72727272",
		505 =>	x"72727272",
		506 =>	x"72727272",
		507 =>	x"397E7F80",
		508 =>	x"81767778",
		509 =>	x"72727272",
		510 =>	x"72727272",
		511 =>	x"82150204", -- IMG_16x16_4intersection
		512 =>	x"8384850D",
		513 =>	x"0D0D0D83",
		514 =>	x"04040282",
		515 =>	x"08020430",
		516 =>	x"860D0D0D",
		517 =>	x"0D0D0D86",
		518 =>	x"87040208",
		519 =>	x"030C0488",
		520 =>	x"0D0D0D0D",
		521 =>	x"0D0D0D0D",
		522 =>	x"0D898A03",
		523 =>	x"1C1C1C8B",
		524 =>	x"0D0D0D0D",
		525 =>	x"0D0D0D0D",
		526 =>	x"0D0D8B1C",
		527 =>	x"84860D85",
		528 =>	x"0D0D0D0D",
		529 =>	x"0D0D0D0D",
		530 =>	x"0D0D0D0D",
		531 =>	x"8C0D0D0D",
		532 =>	x"0D0D0D0D",
		533 =>	x"0D0D0D0D",
		534 =>	x"0D0D0D0D",
		535 =>	x"0D0D0D0D",
		536 =>	x"0D0D0D0D",
		537 =>	x"0D0D0D0D",
		538 =>	x"0D0D0D0D",
		539 =>	x"0D0D0D0D",
		540 =>	x"0D0D0D0D",
		541 =>	x"0D0D0D0D",
		542 =>	x"0D0D0D0D",
		543 =>	x"0D0D0D0D",
		544 =>	x"0D0D0D0D",
		545 =>	x"0D0D0D0D",
		546 =>	x"0D0D0D0D",
		547 =>	x"0D0D0D0D",
		548 =>	x"0D0D0D0D",
		549 =>	x"0D0D0D0D",
		550 =>	x"0D0D0D0D",
		551 =>	x"0D0D0D0D",
		552 =>	x"0D0D0D0D",
		553 =>	x"0D0D0D0D",
		554 =>	x"0D0D0D0D",
		555 =>	x"8D0D0D0D",
		556 =>	x"0D0D0D0D",
		557 =>	x"0D0D0D0D",
		558 =>	x"0D0D0D0D",
		559 =>	x"8E8F0D0D",
		560 =>	x"0D0D0D0D",
		561 =>	x"0D0D0D0D",
		562 =>	x"0D0D908E",
		563 =>	x"2626910D",
		564 =>	x"0D0D0D0D",
		565 =>	x"0D0D0D0D",
		566 =>	x"0D922626",
		567 =>	x"0202041C",
		568 =>	x"930D0D0D",
		569 =>	x"0D0D0D0D",
		570 =>	x"0D040202",
		571 =>	x"82029404",
		572 =>	x"8C0D0D0D",
		573 =>	x"0D0D0D0D",
		574 =>	x"0D040282",
		575 =>	x"82828282", -- IMG_16x16_4middle_horizontal
		576 =>	x"82828282",
		577 =>	x"82828282",
		578 =>	x"82828282",
		579 =>	x"35358282",
		580 =>	x"82353535",
		581 =>	x"35823535",
		582 =>	x"82828235",
		583 =>	x"342D2D34",
		584 =>	x"34343434",
		585 =>	x"2E34342D",
		586 =>	x"342D2D34",
		587 =>	x"04040404",
		588 =>	x"04040404",
		589 =>	x"04040404",
		590 =>	x"042A0404",
		591 =>	x"95108383",
		592 =>	x"10838383",
		593 =>	x"83838396",
		594 =>	x"97839797",
		595 =>	x"83838383",
		596 =>	x"83838383",
		597 =>	x"83838383",
		598 =>	x"83838383",
		599 =>	x"83838383",
		600 =>	x"83838383",
		601 =>	x"83838383",
		602 =>	x"83838383",
		603 =>	x"83838383",
		604 =>	x"83838383",
		605 =>	x"83838383",
		606 =>	x"83838383",
		607 =>	x"83838383",
		608 =>	x"83838383",
		609 =>	x"83838383",
		610 =>	x"83838383",
		611 =>	x"98838383",
		612 =>	x"83838383",
		613 =>	x"83838383",
		614 =>	x"83838383",
		615 =>	x"83838383",
		616 =>	x"83838383",
		617 =>	x"83838383",
		618 =>	x"83838383",
		619 =>	x"83838383",
		620 =>	x"83838383",
		621 =>	x"83838383",
		622 =>	x"83839983",
		623 =>	x"83838383",
		624 =>	x"83838383",
		625 =>	x"83838383",
		626 =>	x"8383049A",
		627 =>	x"9B838383",
		628 =>	x"83839C04",
		629 =>	x"9D838383",
		630 =>	x"839C0404",
		631 =>	x"142D9E14",
		632 =>	x"022D149E",
		633 =>	x"2D9E2D2D",
		634 =>	x"9E2D9E9E",
		635 =>	x"029F9F9F",
		636 =>	x"82829F9F",
		637 =>	x"9F9F9F82",
		638 =>	x"9F828282",
		639 =>	x"36373800", -- IMG_16x16_5end_up
		640 =>	x"393A3B3C",
		641 =>	x"3D3E3F40",
		642 =>	x"00414243",
		643 =>	x"44454647",
		644 =>	x"48493F40",
		645 =>	x"4A4B4C4D",
		646 =>	x"4E4F5000",
		647 =>	x"51525354",
		648 =>	x"55565758",
		649 =>	x"595A5B5C",
		650 =>	x"5D5E5F60",
		651 =>	x"00006162",
		652 =>	x"6364654D",
		653 =>	x"66676800",
		654 =>	x"696A6B39",
		655 =>	x"00000000",
		656 =>	x"00000000",
		657 =>	x"00000000",
		658 =>	x"00000000",
		659 =>	x"00000000",
		660 =>	x"00000000",
		661 =>	x"00000000",
		662 =>	x"00000000",
		663 =>	x"00000000",
		664 =>	x"006C6D6E",
		665 =>	x"6F707100",
		666 =>	x"00000000",
		667 =>	x"00000000",
		668 =>	x"00000000",
		669 =>	x"00000000",
		670 =>	x"00000000",
		671 =>	x"00000000",
		672 =>	x"00000000",
		673 =>	x"00000000",
		674 =>	x"00000000",
		675 =>	x"00000000",
		676 =>	x"00000000",
		677 =>	x"00000000",
		678 =>	x"00000000",
		679 =>	x"00000000",
		680 =>	x"00000000",
		681 =>	x"00000000",
		682 =>	x"00000000",
		683 =>	x"00000000",
		684 =>	x"00000000",
		685 =>	x"00000000",
		686 =>	x"00000000",
		687 =>	x"72727374",
		688 =>	x"75767778",
		689 =>	x"797A7B7C",
		690 =>	x"7D000000",
		691 =>	x"72727272",
		692 =>	x"72727272",
		693 =>	x"72727272",
		694 =>	x"72727272",
		695 =>	x"72727272",
		696 =>	x"72727272",
		697 =>	x"72727272",
		698 =>	x"72727272",
		699 =>	x"397E7F80",
		700 =>	x"81767778",
		701 =>	x"72727272",
		702 =>	x"72727272",
		703 =>	x"82150204", -- IMG_16x16_5intersection
		704 =>	x"17171717",
		705 =>	x"17171704",
		706 =>	x"04028282",
		707 =>	x"82020204",
		708 =>	x"A0171717",
		709 =>	x"17171717",
		710 =>	x"04020282",
		711 =>	x"02020204",
		712 =>	x"17171717",
		713 =>	x"17171717",
		714 =>	x"04030202",
		715 =>	x"A1040404",
		716 =>	x"17171717",
		717 =>	x"17171717",
		718 =>	x"040404A1",
		719 =>	x"04040404",
		720 =>	x"17171717",
		721 =>	x"17171717",
		722 =>	x"04040404",
		723 =>	x"A2A3A3A3",
		724 =>	x"17171717",
		725 =>	x"17171717",
		726 =>	x"A2A3A3A2",
		727 =>	x"A41717A4",
		728 =>	x"A4A51717",
		729 =>	x"17171717",
		730 =>	x"17171717",
		731 =>	x"A6171717",
		732 =>	x"17171717",
		733 =>	x"17171717",
		734 =>	x"17171717",
		735 =>	x"17171717",
		736 =>	x"17171717",
		737 =>	x"17171717",
		738 =>	x"17171717",
		739 =>	x"17171717",
		740 =>	x"17171717",
		741 =>	x"17171717",
		742 =>	x"17171717",
		743 =>	x"A7171717",
		744 =>	x"17171717",
		745 =>	x"171717A8",
		746 =>	x"17171717",
		747 =>	x"13111317",
		748 =>	x"171717A2",
		749 =>	x"17171717",
		750 =>	x"A91717AA",
		751 =>	x"060404A2",
		752 =>	x"17171717",
		753 =>	x"17171717",
		754 =>	x"04060606",
		755 =>	x"020304AB",
		756 =>	x"17171717",
		757 =>	x"17171717",
		758 =>	x"04020202",
		759 =>	x"02020317",
		760 =>	x"17171717",
		761 =>	x"17171704",
		762 =>	x"04020202",
		763 =>	x"82020204",
		764 =>	x"17171717",
		765 =>	x"17171704",
		766 =>	x"26028282",
		767 =>	x"82828282", -- IMG_16x16_5middle_horizontal
		768 =>	x"82828282",
		769 =>	x"82828282",
		770 =>	x"82828282",
		771 =>	x"82828282",
		772 =>	x"82828282",
		773 =>	x"82828282",
		774 =>	x"82828282",
		775 =>	x"02022B02",
		776 =>	x"02020202",
		777 =>	x"02020202",
		778 =>	x"02022B02",
		779 =>	x"2CAC1717",
		780 =>	x"AD170202",
		781 =>	x"2D02022D",
		782 =>	x"0202022D",
		783 =>	x"AEAF1717",
		784 =>	x"1717B02E",
		785 =>	x"04B02D04",
		786 =>	x"2E2D2D04",
		787 =>	x"B1171717",
		788 =>	x"17171717",
		789 =>	x"17171717",
		790 =>	x"17171717",
		791 =>	x"17171717",
		792 =>	x"17171717",
		793 =>	x"17171717",
		794 =>	x"17171717",
		795 =>	x"17171717",
		796 =>	x"17171717",
		797 =>	x"17171717",
		798 =>	x"17171717",
		799 =>	x"17171717",
		800 =>	x"17171717",
		801 =>	x"17171717",
		802 =>	x"17171717",
		803 =>	x"17171717",
		804 =>	x"17171717",
		805 =>	x"17171717",
		806 =>	x"17171717",
		807 =>	x"17171717",
		808 =>	x"17171717",
		809 =>	x"17171717",
		810 =>	x"17171717",
		811 =>	x"A2171717",
		812 =>	x"17171717",
		813 =>	x"17171717",
		814 =>	x"17171717",
		815 =>	x"B2171717",
		816 =>	x"17171717",
		817 =>	x"17171717",
		818 =>	x"17171717",
		819 =>	x"2D2D0202",
		820 =>	x"02020202",
		821 =>	x"02343402",
		822 =>	x"2D020202",
		823 =>	x"02020202",
		824 =>	x"02020202",
		825 =>	x"02020202",
		826 =>	x"02020202",
		827 =>	x"9F828282",
		828 =>	x"82829F82",
		829 =>	x"82828282",
		830 =>	x"82828282",
		831 =>	x"82821A02", -- IMG_16x16_6end_up
		832 =>	x"B3B4B5B5",
		833 =>	x"B5B60602",
		834 =>	x"B7828282",
		835 =>	x"82828202",
		836 =>	x"B3B8B5B5",
		837 =>	x"B5B50602",
		838 =>	x"82828282",
		839 =>	x"82828202",
		840 =>	x"02B6B5B5",
		841 =>	x"B5B50302",
		842 =>	x"82828282",
		843 =>	x"82828202",
		844 =>	x"02B9B5B5",
		845 =>	x"B5B50302",
		846 =>	x"82828282",
		847 =>	x"82828202",
		848 =>	x"BABBB5B5",
		849 =>	x"B5BC0602",
		850 =>	x"82828282",
		851 =>	x"82828202",
		852 =>	x"BDB5B5B5",
		853 =>	x"B5BE0602",
		854 =>	x"82828282",
		855 =>	x"82821A02",
		856 =>	x"BFB5B5B5",
		857 =>	x"B5B50202",
		858 =>	x"82828282",
		859 =>	x"82828202",
		860 =>	x"C0B5B5B5",
		861 =>	x"B5B50302",
		862 =>	x"82828282",
		863 =>	x"82828202",
		864 =>	x"02B5B5B5",
		865 =>	x"B5B5C102",
		866 =>	x"C2828282",
		867 =>	x"82828202",
		868 =>	x"C3B5B5B5",
		869 =>	x"B5C40202",
		870 =>	x"82828282",
		871 =>	x"82828202",
		872 =>	x"C3B6B5B5",
		873 =>	x"B5C50202",
		874 =>	x"82828282",
		875 =>	x"82828202",
		876 =>	x"02B8B5B5",
		877 =>	x"B504C102",
		878 =>	x"C2828282",
		879 =>	x"82828202",
		880 =>	x"B3B6B5B5",
		881 =>	x"B5040302",
		882 =>	x"82828282",
		883 =>	x"82828202",
		884 =>	x"02C6B5B5",
		885 =>	x"B9C70202",
		886 =>	x"82828282",
		887 =>	x"82828282",
		888 =>	x"02B3042E",
		889 =>	x"02020202",
		890 =>	x"82828282",
		891 =>	x"82828282",
		892 =>	x"82020202",
		893 =>	x"0202C882",
		894 =>	x"82828282",
		895 =>	x"82828202", -- IMG_16x16_6intersection
		896 =>	x"0202C9B5",
		897 =>	x"B5B5B602",
		898 =>	x"02828282",
		899 =>	x"82828202",
		900 =>	x"0202B8B5",
		901 =>	x"B5B5B502",
		902 =>	x"02828282",
		903 =>	x"8282821A",
		904 =>	x"0204B5B5",
		905 =>	x"B5B5B502",
		906 =>	x"02828282",
		907 =>	x"82828202",
		908 =>	x"0204B5B5",
		909 =>	x"B5B5B502",
		910 =>	x"02828282",
		911 =>	x"020202B5",
		912 =>	x"B5B5B5B5",
		913 =>	x"B5B5B5B5",
		914 =>	x"B5020202",
		915 =>	x"CA02CBB8",
		916 =>	x"B5B5B5B5",
		917 =>	x"B5B5B5B6",
		918 =>	x"B5B3B304",
		919 =>	x"B8B8B5B5",
		920 =>	x"B5B5B5B5",
		921 =>	x"B5B5B5B5",
		922 =>	x"B5B8B4B8",
		923 =>	x"B5B5B5B5",
		924 =>	x"B5B5B5B5",
		925 =>	x"B5CCB5B5",
		926 =>	x"B5CCB5B5",
		927 =>	x"B5B5B5B5",
		928 =>	x"B5B5B5B5",
		929 =>	x"CCB5B5B5",
		930 =>	x"B5B5B5B5",
		931 =>	x"B5B5B5B5",
		932 =>	x"B5B5B5B5",
		933 =>	x"B5B5B5B5",
		934 =>	x"B5B5B5BC",
		935 =>	x"CDB5B5B5",
		936 =>	x"B5B5B5B5",
		937 =>	x"B5B5B5B5",
		938 =>	x"B5B506C1",
		939 =>	x"02020303",
		940 =>	x"CEB5B5B5",
		941 =>	x"B5B5B5CE",
		942 =>	x"03020202",
		943 =>	x"02020202",
		944 =>	x"0204B5B5",
		945 =>	x"B5B5B502",
		946 =>	x"02020202",
		947 =>	x"82828202",
		948 =>	x"022504B5",
		949 =>	x"B5B5B502",
		950 =>	x"82828282",
		951 =>	x"82828202",
		952 =>	x"020204B5",
		953 =>	x"B5B5B502",
		954 =>	x"02828282",
		955 =>	x"828282CF",
		956 =>	x"020204B5",
		957 =>	x"B5B5B902",
		958 =>	x"02828282",
		959 =>	x"36373800", -- IMG_16x16_6middle_horizontal
		960 =>	x"393A3B3C",
		961 =>	x"3D3E3F40",
		962 =>	x"00414243",
		963 =>	x"44454647",
		964 =>	x"48493F40",
		965 =>	x"4A4B4C4D",
		966 =>	x"4E4F5000",
		967 =>	x"51525354",
		968 =>	x"55565758",
		969 =>	x"595A5B5C",
		970 =>	x"5D5E5F60",
		971 =>	x"00006162",
		972 =>	x"6364654D",
		973 =>	x"66676800",
		974 =>	x"696A6B39",
		975 =>	x"00000000",
		976 =>	x"00000000",
		977 =>	x"00000000",
		978 =>	x"00000000",
		979 =>	x"00000000",
		980 =>	x"00000000",
		981 =>	x"00000000",
		982 =>	x"00000000",
		983 =>	x"00000000",
		984 =>	x"006C6D6E",
		985 =>	x"6F707100",
		986 =>	x"00000000",
		987 =>	x"00000000",
		988 =>	x"00000000",
		989 =>	x"00000000",
		990 =>	x"00000000",
		991 =>	x"00000000",
		992 =>	x"00000000",
		993 =>	x"00000000",
		994 =>	x"00000000",
		995 =>	x"00000000",
		996 =>	x"00000000",
		997 =>	x"00000000",
		998 =>	x"00000000",
		999 =>	x"00000000",
		1000 =>	x"00000000",
		1001 =>	x"00000000",
		1002 =>	x"00000000",
		1003 =>	x"00000000",
		1004 =>	x"00000000",
		1005 =>	x"00000000",
		1006 =>	x"00000000",
		1007 =>	x"72727272",
		1008 =>	x"72727272",
		1009 =>	x"797A7B7C",
		1010 =>	x"7D000000",
		1011 =>	x"72727272",
		1012 =>	x"72727272",
		1013 =>	x"72727272",
		1014 =>	x"72727272",
		1015 =>	x"72727272",
		1016 =>	x"72727272",
		1017 =>	x"72727272",
		1018 =>	x"72727272",
		1019 =>	x"397E7F80",
		1020 =>	x"81767778",
		1021 =>	x"72727272",
		1022 =>	x"72727272",
		1023 =>	x"36373800", -- IMG_16x16_7end_up
		1024 =>	x"393A3B3C",
		1025 =>	x"3D3E3F40",
		1026 =>	x"00414243",
		1027 =>	x"44454647",
		1028 =>	x"48493F40",
		1029 =>	x"4A4B4C4D",
		1030 =>	x"4E4F5000",
		1031 =>	x"51525354",
		1032 =>	x"55565758",
		1033 =>	x"595A5B5C",
		1034 =>	x"5D5E5F60",
		1035 =>	x"00006162",
		1036 =>	x"6364654D",
		1037 =>	x"66676800",
		1038 =>	x"696A6B39",
		1039 =>	x"00000000",
		1040 =>	x"00000000",
		1041 =>	x"00000000",
		1042 =>	x"00000000",
		1043 =>	x"00000000",
		1044 =>	x"00000000",
		1045 =>	x"00000000",
		1046 =>	x"00000000",
		1047 =>	x"00000000",
		1048 =>	x"006C6D6E",
		1049 =>	x"6F707100",
		1050 =>	x"00000000",
		1051 =>	x"00000000",
		1052 =>	x"00000000",
		1053 =>	x"00000000",
		1054 =>	x"00000000",
		1055 =>	x"00000000",
		1056 =>	x"00000000",
		1057 =>	x"00000000",
		1058 =>	x"00000000",
		1059 =>	x"00000000",
		1060 =>	x"00000000",
		1061 =>	x"00000000",
		1062 =>	x"00000000",
		1063 =>	x"00000000",
		1064 =>	x"00000000",
		1065 =>	x"00000000",
		1066 =>	x"00000000",
		1067 =>	x"00000000",
		1068 =>	x"00000000",
		1069 =>	x"00000000",
		1070 =>	x"00000000",
		1071 =>	x"72727374",
		1072 =>	x"75767778",
		1073 =>	x"797A7B7C",
		1074 =>	x"7D000000",
		1075 =>	x"72727272",
		1076 =>	x"72727272",
		1077 =>	x"72727272",
		1078 =>	x"72727272",
		1079 =>	x"72727272",
		1080 =>	x"72727272",
		1081 =>	x"72727272",
		1082 =>	x"72727272",
		1083 =>	x"397E7F80",
		1084 =>	x"81767778",
		1085 =>	x"72727272",
		1086 =>	x"72727272",
		1087 =>	x"82828282", -- IMG_16x16_7middle_horizontal
		1088 =>	x"82828282",
		1089 =>	x"82828282",
		1090 =>	x"82828282",
		1091 =>	x"82828282",
		1092 =>	x"82828282",
		1093 =>	x"82828282",
		1094 =>	x"82828282",
		1095 =>	x"82828282",
		1096 =>	x"82828282",
		1097 =>	x"82828282",
		1098 =>	x"82828282",
		1099 =>	x"82828282",
		1100 =>	x"82828282",
		1101 =>	x"82828282",
		1102 =>	x"82828282",
		1103 =>	x"02028202",
		1104 =>	x"02820282",
		1105 =>	x"82828282",
		1106 =>	x"82828282",
		1107 =>	x"02020202",
		1108 =>	x"02020202",
		1109 =>	x"D0020202",
		1110 =>	x"D002D002",
		1111 =>	x"D1D2D2D2",
		1112 =>	x"D2D2D2D3",
		1113 =>	x"D4D5D6D2",
		1114 =>	x"D2D2D2D6",
		1115 =>	x"D2D2D2D2",
		1116 =>	x"D2D2D2D2",
		1117 =>	x"D2D2D2D2",
		1118 =>	x"D2D2D2D2",
		1119 =>	x"D2D2D2D2",
		1120 =>	x"D2D2D2D2",
		1121 =>	x"D2D2D2D2",
		1122 =>	x"D2D2D2D2",
		1123 =>	x"D2D2D2D2",
		1124 =>	x"D2D2D2D2",
		1125 =>	x"D2D2D2D2",
		1126 =>	x"D2D2D2D2",
		1127 =>	x"02020202",
		1128 =>	x"02020202",
		1129 =>	x"02D70202",
		1130 =>	x"02020202",
		1131 =>	x"82028202",
		1132 =>	x"82028202",
		1133 =>	x"D8D80202",
		1134 =>	x"82028282",
		1135 =>	x"82828282",
		1136 =>	x"82828282",
		1137 =>	x"82828282",
		1138 =>	x"82828282",
		1139 =>	x"82828282",
		1140 =>	x"82828282",
		1141 =>	x"82828282",
		1142 =>	x"82828282",
		1143 =>	x"82828282",
		1144 =>	x"82828282",
		1145 =>	x"82828282",
		1146 =>	x"82828282",
		1147 =>	x"82828282",
		1148 =>	x"82828282",
		1149 =>	x"82828282",
		1150 =>	x"82828282",
		1151 =>	x"01010101", -- IMG_16x16_background
		1152 =>	x"01010101",
		1153 =>	x"01010101",
		1154 =>	x"01010101",
		1155 =>	x"01010101",
		1156 =>	x"01010101",
		1157 =>	x"01010101",
		1158 =>	x"01010101",
		1159 =>	x"01010101",
		1160 =>	x"01010101",
		1161 =>	x"01010101",
		1162 =>	x"01010101",
		1163 =>	x"01010101",
		1164 =>	x"01010101",
		1165 =>	x"01010101",
		1166 =>	x"01010101",
		1167 =>	x"01010101",
		1168 =>	x"01010101",
		1169 =>	x"01010101",
		1170 =>	x"01010101",
		1171 =>	x"01010101",
		1172 =>	x"01010101",
		1173 =>	x"01010101",
		1174 =>	x"01010101",
		1175 =>	x"01010101",
		1176 =>	x"01010101",
		1177 =>	x"01010101",
		1178 =>	x"01010101",
		1179 =>	x"01010101",
		1180 =>	x"01010101",
		1181 =>	x"01010101",
		1182 =>	x"01010101",
		1183 =>	x"01010101",
		1184 =>	x"01010101",
		1185 =>	x"01010101",
		1186 =>	x"01010101",
		1187 =>	x"01010101",
		1188 =>	x"01010101",
		1189 =>	x"01010101",
		1190 =>	x"01010101",
		1191 =>	x"01010101",
		1192 =>	x"01010101",
		1193 =>	x"01010101",
		1194 =>	x"01010101",
		1195 =>	x"01010101",
		1196 =>	x"01010101",
		1197 =>	x"01010101",
		1198 =>	x"01010101",
		1199 =>	x"01010101",
		1200 =>	x"01010101",
		1201 =>	x"01010101",
		1202 =>	x"01010101",
		1203 =>	x"01010101",
		1204 =>	x"01010101",
		1205 =>	x"01010101",
		1206 =>	x"01010101",
		1207 =>	x"01010101",
		1208 =>	x"01010101",
		1209 =>	x"01010101",
		1210 =>	x"01010101",
		1211 =>	x"01010101",
		1212 =>	x"01010101",
		1213 =>	x"01010101",
		1214 =>	x"01010101",
		1215 =>	x"82828282", -- IMG_16x16_block
		1216 =>	x"82828282",
		1217 =>	x"82828282",
		1218 =>	x"8282D901",
		1219 =>	x"DADADADA",
		1220 =>	x"DADADADA",
		1221 =>	x"DADADADA",
		1222 =>	x"DADAD901",
		1223 =>	x"DADADADA",
		1224 =>	x"DADADADA",
		1225 =>	x"DADADADA",
		1226 =>	x"DADAD901",
		1227 =>	x"DADADADA",
		1228 =>	x"DADADADA",
		1229 =>	x"DADADADA",
		1230 =>	x"DADAD901",
		1231 =>	x"DADADADA",
		1232 =>	x"DADADADA",
		1233 =>	x"DADADADA",
		1234 =>	x"DADAD901",
		1235 =>	x"DADADADA",
		1236 =>	x"DADADADA",
		1237 =>	x"DADADADA",
		1238 =>	x"DADAD901",
		1239 =>	x"DADADADA",
		1240 =>	x"DADADADA",
		1241 =>	x"DADADADA",
		1242 =>	x"DADAD901",
		1243 =>	x"DADADADA",
		1244 =>	x"DADADADA",
		1245 =>	x"DADADADA",
		1246 =>	x"DADAD901",
		1247 =>	x"DADADADA",
		1248 =>	x"DADADADA",
		1249 =>	x"DADADADA",
		1250 =>	x"DADAD901",
		1251 =>	x"DADADADA",
		1252 =>	x"DADADADA",
		1253 =>	x"DADADADA",
		1254 =>	x"DADAD901",
		1255 =>	x"DADADADA",
		1256 =>	x"DADADADA",
		1257 =>	x"DADADADA",
		1258 =>	x"DADAD901",
		1259 =>	x"DADADADA",
		1260 =>	x"DADADADA",
		1261 =>	x"DADADADA",
		1262 =>	x"DADAD901",
		1263 =>	x"DADADADA",
		1264 =>	x"DADADADA",
		1265 =>	x"DADADADA",
		1266 =>	x"DADAD901",
		1267 =>	x"DADADADA",
		1268 =>	x"DADADADA",
		1269 =>	x"DADADADA",
		1270 =>	x"DADAD901",
		1271 =>	x"D9D9D9D9",
		1272 =>	x"D9D9D9D9",
		1273 =>	x"D9D9D9D9",
		1274 =>	x"D9DAD901",
		1275 =>	x"D9D9D9D9",
		1276 =>	x"D9D9D9D9",
		1277 =>	x"D9D9D9D9",
		1278 =>	x"D9D9D901",
		1279 =>	x"01010101", -- IMG_16x16_bomb
		1280 =>	x"01010101",
		1281 =>	x"01010101",
		1282 =>	x"01010101",
		1283 =>	x"01010101",
		1284 =>	x"01010101",
		1285 =>	x"01828282",
		1286 =>	x"01820182",
		1287 =>	x"01010101",
		1288 =>	x"01D9D9D9",
		1289 =>	x"8282D9D9",
		1290 =>	x"01010101",
		1291 =>	x"010101D9",
		1292 =>	x"D9D9D9D9",
		1293 =>	x"82D9D9D9",
		1294 =>	x"D9018201",
		1295 =>	x"0101D9D9",
		1296 =>	x"8282D9D9",
		1297 =>	x"82D9D9D9",
		1298 =>	x"D9D90101",
		1299 =>	x"01D9D982",
		1300 =>	x"82D9D9D9",
		1301 =>	x"D9D9D9D9",
		1302 =>	x"D9D9D901",
		1303 =>	x"01D9D982",
		1304 =>	x"82D9D9D9",
		1305 =>	x"D9D9D9D9",
		1306 =>	x"D9D9D901",
		1307 =>	x"D9D98282",
		1308 =>	x"D9D9D9D9",
		1309 =>	x"D9D9D9D9",
		1310 =>	x"D9D9D9D9",
		1311 =>	x"D9D98282",
		1312 =>	x"D9D9D9D9",
		1313 =>	x"D9D9D9D9",
		1314 =>	x"D9D9D9D9",
		1315 =>	x"D9D9D9D9",
		1316 =>	x"D9D9D9D9",
		1317 =>	x"D9D9D9D9",
		1318 =>	x"D9D9D9D9",
		1319 =>	x"D9D9D9D9",
		1320 =>	x"D9D9D9D9",
		1321 =>	x"D9D9D9D9",
		1322 =>	x"D9D9D9D9",
		1323 =>	x"D9D9D9D9",
		1324 =>	x"D9D9D9D9",
		1325 =>	x"D9D9D9D9",
		1326 =>	x"D9D9D9D9",
		1327 =>	x"01D9D9D9",
		1328 =>	x"D9D9D9D9",
		1329 =>	x"D9D9D9D9",
		1330 =>	x"D9D9D901",
		1331 =>	x"01D9D9D9",
		1332 =>	x"D9D9D9D9",
		1333 =>	x"D9D9D9D9",
		1334 =>	x"D9D9D901",
		1335 =>	x"0101D9D9",
		1336 =>	x"D9D9D9D9",
		1337 =>	x"D9D9D9D9",
		1338 =>	x"D9D90101",
		1339 =>	x"010101D9",
		1340 =>	x"D9D9D9D9",
		1341 =>	x"D9D9D9D9",
		1342 =>	x"D9010101",
		1343 =>	x"01010101", -- IMG_16x16_bomberman
		1344 =>	x"01828282",
		1345 =>	x"82828201",
		1346 =>	x"01010101",
		1347 =>	x"01010101",
		1348 =>	x"82828282",
		1349 =>	x"82828282",
		1350 =>	x"01010101",
		1351 =>	x"01010101",
		1352 =>	x"82DB01DB",
		1353 =>	x"DB01DB82",
		1354 =>	x"01010101",
		1355 =>	x"01010101",
		1356 =>	x"82DB01DB",
		1357 =>	x"DB01DB82",
		1358 =>	x"01010101",
		1359 =>	x"01010101",
		1360 =>	x"82828282",
		1361 =>	x"82828282",
		1362 =>	x"01010101",
		1363 =>	x"01010101",
		1364 =>	x"01828282",
		1365 =>	x"82828201",
		1366 =>	x"01010101",
		1367 =>	x"01010101",
		1368 =>	x"0101DCDC",
		1369 =>	x"DCDC0101",
		1370 =>	x"01010101",
		1371 =>	x"01010101",
		1372 =>	x"8282DCDC",
		1373 =>	x"DCDC8282",
		1374 =>	x"01010101",
		1375 =>	x"01010182",
		1376 =>	x"82DCDCDC",
		1377 =>	x"DCDCDC82",
		1378 =>	x"82010101",
		1379 =>	x"0101DBDB",
		1380 =>	x"82DCDCDC",
		1381 =>	x"DCDCDC82",
		1382 =>	x"DBDB0101",
		1383 =>	x"0101DBDB",
		1384 =>	x"01DCDCDC",
		1385 =>	x"DCDCDC01",
		1386 =>	x"DBDB0101",
		1387 =>	x"01010101",
		1388 =>	x"01DCDCDC",
		1389 =>	x"DCDCDC01",
		1390 =>	x"01010101",
		1391 =>	x"01010101",
		1392 =>	x"018282DC",
		1393 =>	x"DC828201",
		1394 =>	x"01010101",
		1395 =>	x"01010101",
		1396 =>	x"01828201",
		1397 =>	x"01828201",
		1398 =>	x"01010101",
		1399 =>	x"01010101",
		1400 =>	x"01DBDB01",
		1401 =>	x"01DBDB01",
		1402 =>	x"01010101",
		1403 =>	x"01010101",
		1404 =>	x"01DBDB01",
		1405 =>	x"01DBDB01",
		1406 =>	x"01010101",
		1407 =>	x"01010101", -- IMG_16x16_bomberman_bomb
		1408 =>	x"01828282",
		1409 =>	x"82828201",
		1410 =>	x"01010101",
		1411 =>	x"01010101",
		1412 =>	x"82828282",
		1413 =>	x"82828282",
		1414 =>	x"01010101",
		1415 =>	x"01010101",
		1416 =>	x"82DB01DB",
		1417 =>	x"DB01DB82",
		1418 =>	x"01010101",
		1419 =>	x"01010100",
		1420 =>	x"82DB01DB",
		1421 =>	x"DB01DB82",
		1422 =>	x"00010101",
		1423 =>	x"01010000",
		1424 =>	x"82828282",
		1425 =>	x"82828282",
		1426 =>	x"00000101",
		1427 =>	x"01000000",
		1428 =>	x"00828282",
		1429 =>	x"82828200",
		1430 =>	x"00000001",
		1431 =>	x"01000000",
		1432 =>	x"0000DCDC",
		1433 =>	x"DCDC0000",
		1434 =>	x"00000001",
		1435 =>	x"00000000",
		1436 =>	x"8282DCDC",
		1437 =>	x"DCDC8282",
		1438 =>	x"00000000",
		1439 =>	x"00000082",
		1440 =>	x"82DCDCDC",
		1441 =>	x"DCDCDC82",
		1442 =>	x"82000000",
		1443 =>	x"0000DBDB",
		1444 =>	x"82DCDCDC",
		1445 =>	x"DCDCDC82",
		1446 =>	x"DBDB0000",
		1447 =>	x"0000DBDB",
		1448 =>	x"00DCDCDC",
		1449 =>	x"DCDCDC00",
		1450 =>	x"DBDB0000",
		1451 =>	x"00000000",
		1452 =>	x"00DCDCDC",
		1453 =>	x"DCDCDC00",
		1454 =>	x"00000000",
		1455 =>	x"01000000",
		1456 =>	x"008282DC",
		1457 =>	x"DC828200",
		1458 =>	x"00000001",
		1459 =>	x"01000000",
		1460 =>	x"00828200",
		1461 =>	x"00828200",
		1462 =>	x"00000001",
		1463 =>	x"01010000",
		1464 =>	x"00DBDB00",
		1465 =>	x"00DBDB00",
		1466 =>	x"00000101",
		1467 =>	x"01010100",
		1468 =>	x"00DBDB00",
		1469 =>	x"00DBDB00",
		1470 =>	x"00010101",
		1471 =>	x"D9D9D9D9", -- IMG_16x16_brick
		1472 =>	x"D9D9D9D9",
		1473 =>	x"D9D9D9D9",
		1474 =>	x"D9D9D9D9",
		1475 =>	x"D9828282",
		1476 =>	x"82828282",
		1477 =>	x"82828282",
		1478 =>	x"828282D9",
		1479 =>	x"82DADADA",
		1480 =>	x"DADADADA",
		1481 =>	x"DADADADA",
		1482 =>	x"DADADAD9",
		1483 =>	x"82DADADA",
		1484 =>	x"DADADADA",
		1485 =>	x"DADADADA",
		1486 =>	x"DADADAD9",
		1487 =>	x"82DADADA",
		1488 =>	x"DADADADA",
		1489 =>	x"DADADADA",
		1490 =>	x"DADADAD9",
		1491 =>	x"D9D9D9D9",
		1492 =>	x"D9D9D9D9",
		1493 =>	x"D9D9D9D9",
		1494 =>	x"D9D9D9D9",
		1495 =>	x"82828282",
		1496 =>	x"82D9D982",
		1497 =>	x"82828282",
		1498 =>	x"82828282",
		1499 =>	x"DADADADA",
		1500 =>	x"DAD982DA",
		1501 =>	x"DADADADA",
		1502 =>	x"DADADADA",
		1503 =>	x"DADADADA",
		1504 =>	x"DAD982DA",
		1505 =>	x"DADADADA",
		1506 =>	x"DADADADA",
		1507 =>	x"DADADADA",
		1508 =>	x"DAD982DA",
		1509 =>	x"DADADADA",
		1510 =>	x"DADADADA",
		1511 =>	x"D9D9D9D9",
		1512 =>	x"D9D9D9D9",
		1513 =>	x"D9D9D9D9",
		1514 =>	x"D9D9D9D9",
		1515 =>	x"82828282",
		1516 =>	x"82828282",
		1517 =>	x"82D9D982",
		1518 =>	x"82828282",
		1519 =>	x"DADADADA",
		1520 =>	x"DADADADA",
		1521 =>	x"DAD982DA",
		1522 =>	x"DADADADA",
		1523 =>	x"DADADADA",
		1524 =>	x"DADADADA",
		1525 =>	x"DAD982DA",
		1526 =>	x"DADADADA",
		1527 =>	x"DADADADA",
		1528 =>	x"DADADADA",
		1529 =>	x"DAD982DA",
		1530 =>	x"DADADADA",
		1531 =>	x"D9D9D9D9",
		1532 =>	x"D9D9D9D9",
		1533 =>	x"D9D9D9D9",
		1534 =>	x"D9D9D9D9",
		1535 =>	x"D9DDDDDD", -- IMG_16x16_door
		1536 =>	x"DDDDD9DD",
		1537 =>	x"DDDDDDDD",
		1538 =>	x"D9D90101",
		1539 =>	x"DDDDDEDE",
		1540 =>	x"DEDDD9DD",
		1541 =>	x"DEDEDEDD",
		1542 =>	x"DDD90101",
		1543 =>	x"DDDEDEDD",
		1544 =>	x"DEDDD9DD",
		1545 =>	x"DEDDDEDE",
		1546 =>	x"DDDD0101",
		1547 =>	x"DDDEDEDE",
		1548 =>	x"DEDDD9DD",
		1549 =>	x"DEDEDEDE",
		1550 =>	x"DDDD0101",
		1551 =>	x"DDDEDEDE",
		1552 =>	x"DEDDD9DD",
		1553 =>	x"DEDEDEDE",
		1554 =>	x"DDD90101",
		1555 =>	x"DDDEDED9",
		1556 =>	x"DEDDD9DD",
		1557 =>	x"DED9DEDE",
		1558 =>	x"DDD90101",
		1559 =>	x"DDDEDDD9",
		1560 =>	x"DDDDDDDD",
		1561 =>	x"DDD9DDDE",
		1562 =>	x"DDD90101",
		1563 =>	x"DDDEDDD9",
		1564 =>	x"DDDDDDDD",
		1565 =>	x"DDD9DDDE",
		1566 =>	x"DDD90101",
		1567 =>	x"DDDEDED9",
		1568 =>	x"DEDDD9DD",
		1569 =>	x"DED9DEDE",
		1570 =>	x"DDD90101",
		1571 =>	x"DDDEDEDE",
		1572 =>	x"DEDDD9DD",
		1573 =>	x"DEDEDEDE",
		1574 =>	x"DDD90101",
		1575 =>	x"DDDEDEDE",
		1576 =>	x"DEDDD9DD",
		1577 =>	x"DEDEDEDE",
		1578 =>	x"DDDD0101",
		1579 =>	x"DDDEDEDD",
		1580 =>	x"DEDDD9DD",
		1581 =>	x"DEDDDEDE",
		1582 =>	x"DDDD0101",
		1583 =>	x"DDDDDEDE",
		1584 =>	x"DEDDD9DD",
		1585 =>	x"DEDEDEDD",
		1586 =>	x"DDD90101",
		1587 =>	x"D9DDDDDD",
		1588 =>	x"DDDDD9DD",
		1589 =>	x"DDDDDDDD",
		1590 =>	x"D9D90101",
		1591 =>	x"01010101",
		1592 =>	x"01010101",
		1593 =>	x"01010101",
		1594 =>	x"01010101",
		1595 =>	x"01010101",
		1596 =>	x"01010101",
		1597 =>	x"01010101",
		1598 =>	x"01010101",
		1599 =>	x"01010101", -- IMG_16x16_enemy
		1600 =>	x"01010101",
		1601 =>	x"01010101",
		1602 =>	x"01010101",
		1603 =>	x"01010101",
		1604 =>	x"01010101",
		1605 =>	x"01010101",
		1606 =>	x"01010101",
		1607 =>	x"01010101",
		1608 =>	x"D9D9D9D9",
		1609 =>	x"D9D9D9D9",
		1610 =>	x"01010101",
		1611 =>	x"0101D9D9",
		1612 =>	x"D9DBDBDB",
		1613 =>	x"DBDBDBD9",
		1614 =>	x"D9D90101",
		1615 =>	x"01D9D9DB",
		1616 =>	x"DBDBDBDB",
		1617 =>	x"DBDBDBDB",
		1618 =>	x"DBD9D901",
		1619 =>	x"D9D9DBDB",
		1620 =>	x"DBDBDBDB",
		1621 =>	x"DBDBDBDB",
		1622 =>	x"DBDBD9D9",
		1623 =>	x"D9DBDBDB",
		1624 =>	x"DB8282DB",
		1625 =>	x"DB8282DB",
		1626 =>	x"DBDBDBD9",
		1627 =>	x"D9DBDBDB",
		1628 =>	x"DBD982DB",
		1629 =>	x"DBD982DB",
		1630 =>	x"DBDBDBD9",
		1631 =>	x"D9DBDBDB",
		1632 =>	x"DBD982DB",
		1633 =>	x"DBD982DB",
		1634 =>	x"DBDBDBD9",
		1635 =>	x"D9D9DBDB",
		1636 =>	x"DBDBDBDB",
		1637 =>	x"DBDBDBDB",
		1638 =>	x"DBDBD9D9",
		1639 =>	x"01D9DBDB",
		1640 =>	x"DBDBDBDB",
		1641 =>	x"DBDBDBDB",
		1642 =>	x"DBDBD901",
		1643 =>	x"01D9D9DB",
		1644 =>	x"DBDBDBD9",
		1645 =>	x"D9DBDBDB",
		1646 =>	x"DBD9D901",
		1647 =>	x"0101D9D9",
		1648 =>	x"D9DBDBDB",
		1649 =>	x"DBDBDBD9",
		1650 =>	x"D9D90101",
		1651 =>	x"01010101",
		1652 =>	x"D9D9D9DB",
		1653 =>	x"DBD9D9D9",
		1654 =>	x"01010101",
		1655 =>	x"01010101",
		1656 =>	x"0101D982",
		1657 =>	x"82D90101",
		1658 =>	x"01010101",
		1659 =>	x"01010101",
		1660 =>	x"0101D9D9",
		1661 =>	x"D9D90101",
		1662 =>	x"01010101",
		1663 =>	x"02020202", -- IMG_16x16_plus_bomb
		1664 =>	x"02020202",
		1665 =>	x"02020202",
		1666 =>	x"02020202",
		1667 =>	x"02121212",
		1668 =>	x"12121212",
		1669 =>	x"12828282",
		1670 =>	x"12121202",
		1671 =>	x"02121212",
		1672 =>	x"12D9D9D9",
		1673 =>	x"8282D9D9",
		1674 =>	x"12121202",
		1675 =>	x"021212D9",
		1676 =>	x"D9D9D9D9",
		1677 =>	x"82D9D9D9",
		1678 =>	x"D9121202",
		1679 =>	x"0212D9D9",
		1680 =>	x"8282D9D9",
		1681 =>	x"82D9D9D9",
		1682 =>	x"D9D91202",
		1683 =>	x"02D9D982",
		1684 =>	x"82D9D9D9",
		1685 =>	x"D9D9D9D9",
		1686 =>	x"D9D9D902",
		1687 =>	x"02D9D982",
		1688 =>	x"82D9D9D9",
		1689 =>	x"D9D9D9D9",
		1690 =>	x"D9D9D902",
		1691 =>	x"02D98282",
		1692 =>	x"D9D9D9D9",
		1693 =>	x"D9D9D9D9",
		1694 =>	x"D9D9D902",
		1695 =>	x"02D98282",
		1696 =>	x"D9D9D9D9",
		1697 =>	x"D9D9D9D9",
		1698 =>	x"D9D9D902",
		1699 =>	x"02D9D9D9",
		1700 =>	x"D9D9D9D9",
		1701 =>	x"D9D9D9D9",
		1702 =>	x"D9D9D902",
		1703 =>	x"02D9D9D9",
		1704 =>	x"D9D9D9D9",
		1705 =>	x"D9D9D9D9",
		1706 =>	x"D9D9D902",
		1707 =>	x"02D9D9D9",
		1708 =>	x"D9D9D9D9",
		1709 =>	x"D9D9D9D9",
		1710 =>	x"D9D9D902",
		1711 =>	x"02D9D9D9",
		1712 =>	x"D9D9D9D9",
		1713 =>	x"D9D9D9D9",
		1714 =>	x"D9D9D902",
		1715 =>	x"02D9D9D9",
		1716 =>	x"D9D9D9D9",
		1717 =>	x"D9D9D9D9",
		1718 =>	x"D9D9D902",
		1719 =>	x"0212D9D9",
		1720 =>	x"D9D9D9D9",
		1721 =>	x"D9D9D9D9",
		1722 =>	x"D9D91202",
		1723 =>	x"02020202",
		1724 =>	x"02020202",
		1725 =>	x"02020202",
		1726 =>	x"02020202",
		1727 =>	x"DFDFDFDF", -- IMG_16x16_plus_explosion
		1728 =>	x"DFDFDFDF",
		1729 =>	x"DFDFDFDF",
		1730 =>	x"DFDFDFDF",
		1731 =>	x"DF121212",
		1732 =>	x"12121212",
		1733 =>	x"12121212",
		1734 =>	x"121212DF",
		1735 =>	x"DF121212",
		1736 =>	x"12121202",
		1737 =>	x"02121212",
		1738 =>	x"121212DF",
		1739 =>	x"DF121212",
		1740 =>	x"12121202",
		1741 =>	x"02121212",
		1742 =>	x"121212DF",
		1743 =>	x"DF121212",
		1744 =>	x"1212022E",
		1745 =>	x"2E021212",
		1746 =>	x"121212DF",
		1747 =>	x"DF121212",
		1748 =>	x"1202022E",
		1749 =>	x"2E020212",
		1750 =>	x"121212DF",
		1751 =>	x"DF121212",
		1752 =>	x"02022E12",
		1753 =>	x"122E0202",
		1754 =>	x"121212DF",
		1755 =>	x"DF120202",
		1756 =>	x"2E2E1212",
		1757 =>	x"12122E2E",
		1758 =>	x"020212DF",
		1759 =>	x"DF120202",
		1760 =>	x"2E2E1212",
		1761 =>	x"12122E2E",
		1762 =>	x"020212DF",
		1763 =>	x"DF121212",
		1764 =>	x"02022E12",
		1765 =>	x"122E0202",
		1766 =>	x"121212DF",
		1767 =>	x"DF121212",
		1768 =>	x"1202022E",
		1769 =>	x"2E020212",
		1770 =>	x"121212DF",
		1771 =>	x"DF121212",
		1772 =>	x"1212022E",
		1773 =>	x"2E021212",
		1774 =>	x"121212DF",
		1775 =>	x"DF121212",
		1776 =>	x"12121202",
		1777 =>	x"02121212",
		1778 =>	x"121212DF",
		1779 =>	x"DF121212",
		1780 =>	x"12121202",
		1781 =>	x"02121212",
		1782 =>	x"121212DF",
		1783 =>	x"DF121212",
		1784 =>	x"12121212",
		1785 =>	x"12121212",
		1786 =>	x"121212DF",
		1787 =>	x"DFDFDFDF",
		1788 =>	x"DFDFDFDF",
		1789 =>	x"DFDFDFDF",
		1790 =>	x"DFDFDFDF",


--			***** MAP *****


		1791 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1792 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1793 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1794 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1795 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1796 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1797 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1798 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1799 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1800 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1801 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1802 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1803 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1804 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1805 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1806 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1807 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1808 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1809 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1810 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1811 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1812 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1813 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1814 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1815 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1816 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1817 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1818 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1819 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1820 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1821 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1822 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1823 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1824 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1825 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1826 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1827 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1828 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1829 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1830 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1831 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1832 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1833 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1834 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1835 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1836 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1837 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1838 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1839 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1840 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1841 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1842 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1843 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1844 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1845 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1846 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1847 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1848 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1849 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1850 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1851 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1852 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1853 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1854 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1855 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1856 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1857 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1858 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1859 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1860 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1861 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1862 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1863 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1864 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1865 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1866 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1867 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1868 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1869 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1870 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1871 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1872 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1873 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1874 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1875 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1876 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1877 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1878 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1879 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1880 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1881 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1882 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1883 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1884 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1885 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1886 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1887 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1888 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1889 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1890 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1891 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1892 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1893 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1894 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1895 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1896 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1897 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1898 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1899 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1900 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1901 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1902 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1903 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1904 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1905 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1906 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1907 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1908 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1909 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1910 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1911 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1912 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1913 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1914 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1915 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1916 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1917 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1918 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1919 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1920 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1921 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1922 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1923 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1924 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1925 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1926 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1927 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1928 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1929 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1930 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1931 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1932 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1933 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1934 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1935 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1936 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1937 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1938 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1939 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1940 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1941 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1942 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1943 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1944 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1945 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1946 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1947 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1948 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1949 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1950 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1951 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1952 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1953 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1954 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1955 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1956 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1957 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1958 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1959 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1960 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1961 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1962 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1963 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1964 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1965 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1966 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1967 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1968 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1969 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1970 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1971 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1972 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1973 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1974 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1975 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1976 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1977 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1978 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1979 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1980 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1981 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1982 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1983 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1984 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1985 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1986 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1987 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1988 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1989 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1990 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1991 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1992 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1993 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1994 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1995 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1996 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		1997 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1998 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		1999 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2000 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2001 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2002 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2003 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2004 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2005 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2006 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2007 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2008 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2009 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2010 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2011 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2012 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2013 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2014 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2015 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2016 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2017 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2018 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2019 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2020 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2021 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2022 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2023 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2024 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2025 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2026 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2027 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2028 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2029 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2030 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2031 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2032 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2033 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2034 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2035 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2036 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2037 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2038 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2039 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2040 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2041 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2042 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2043 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2044 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2045 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2046 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2047 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2048 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2049 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2050 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2051 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2052 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2053 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2054 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2055 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2056 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2057 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2058 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2059 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2060 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2061 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2062 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2063 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2064 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2065 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2066 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2067 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2068 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2069 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2070 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2071 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2072 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2073 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2074 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2075 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2076 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2077 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2078 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2079 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2080 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2081 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2082 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2083 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2084 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2085 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2086 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2087 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2088 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2089 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2090 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2091 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2092 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2093 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2094 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2095 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2096 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2097 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2098 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2099 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2100 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2101 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2102 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2103 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2104 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2105 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2106 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2107 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2108 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2109 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2110 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2111 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2112 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2113 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2114 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2115 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2116 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2117 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2118 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2119 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2120 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2121 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2122 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2123 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2124 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2125 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2126 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2127 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2128 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2129 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2130 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2131 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2132 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2133 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2134 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2135 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2136 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2137 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2138 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2139 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2140 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2141 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2142 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2143 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2144 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2145 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2146 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2147 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2148 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2149 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2150 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2151 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2152 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2153 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2154 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2155 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2156 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2157 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2158 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2159 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2160 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2161 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2162 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2163 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2164 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2165 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2166 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2167 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2168 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2169 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2170 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2171 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2172 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2173 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2174 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2175 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2176 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2177 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2178 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2179 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2180 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2181 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2182 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2183 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2184 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2185 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2186 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2187 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2188 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2189 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2190 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2191 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2192 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2193 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2194 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2195 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2196 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2197 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2198 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2199 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2200 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2201 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2202 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2203 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2204 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2205 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2206 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2207 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2208 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2209 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2210 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2211 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2212 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2213 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2214 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2215 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2216 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2217 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2218 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2219 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2220 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2221 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2222 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2223 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2224 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2225 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2226 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2227 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2228 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2229 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2230 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2231 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2232 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2233 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2234 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2235 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2236 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2237 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2238 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2239 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2240 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2241 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2242 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2243 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2244 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2245 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2246 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2247 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2248 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2249 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2250 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2251 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2252 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2253 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2254 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2255 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2256 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2257 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2258 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2259 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2260 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2261 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2262 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2263 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2264 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2265 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2266 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2267 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2268 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2269 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2270 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2271 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2272 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2273 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2274 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2275 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2276 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2277 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2278 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2279 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2280 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2281 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2282 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2283 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2284 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2285 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2286 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2287 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2288 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2289 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2290 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2291 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2292 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2293 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2294 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2295 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2296 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2297 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2298 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2299 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2300 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2301 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2302 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2303 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2304 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2305 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2306 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2307 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2308 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2309 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2310 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2311 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2312 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2313 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2314 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2315 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2316 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2317 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2318 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2319 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2320 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2321 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2322 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2323 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2324 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2325 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2326 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2327 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2328 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2329 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2330 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2331 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2332 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2333 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2334 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2335 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2336 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2337 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2338 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2339 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2340 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2341 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2342 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2343 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2344 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2345 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2346 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2347 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2348 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2349 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2350 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2351 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2352 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2353 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2354 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2355 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2356 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2357 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2358 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2359 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2360 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2361 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2362 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2363 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2364 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2365 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2366 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2367 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2368 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2369 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2370 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2371 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2372 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2373 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2374 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2375 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2376 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2377 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2378 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2379 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2380 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2381 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2382 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2383 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2384 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2385 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2386 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2387 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2388 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2389 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2390 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2391 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2392 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2393 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2394 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2395 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2396 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2397 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2398 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2399 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2400 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2401 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2402 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2403 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2404 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2405 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2406 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2407 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2408 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2409 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2410 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2411 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2412 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2413 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2414 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2415 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2416 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2417 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2418 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2419 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2420 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2421 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2422 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2423 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2424 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2425 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2426 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2427 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2428 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2429 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2430 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2431 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2432 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2433 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2434 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2435 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2436 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2437 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2438 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2439 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2440 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2441 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2442 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2443 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2444 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2445 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2446 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2447 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2448 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2449 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2450 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2451 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2452 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2453 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2454 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2455 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2456 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2457 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2458 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2459 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2460 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2461 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2462 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2463 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2464 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2465 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2466 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2467 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2468 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2469 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2470 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2471 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2472 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2473 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2474 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2475 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2476 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2477 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2478 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2479 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2480 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2481 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2482 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2483 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2484 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2485 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2486 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2487 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2488 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2489 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2490 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2491 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2492 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2493 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2494 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2495 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2496 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2497 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2498 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2499 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2500 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2501 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2502 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2503 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2504 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2505 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2506 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2507 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2508 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2509 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2510 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2511 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2512 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2513 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2514 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2515 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2516 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2517 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2518 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2519 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2520 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2521 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2522 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2523 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2524 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2525 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2526 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2527 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2528 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2529 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2530 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2531 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2532 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2533 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2534 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2535 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2536 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2537 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2538 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2539 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2540 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2541 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2542 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2543 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2544 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2545 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2546 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2547 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2548 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2549 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2550 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2551 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2552 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2553 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2554 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2555 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2556 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2557 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2558 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2559 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2560 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2561 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2562 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2563 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2564 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2565 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2566 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2567 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2568 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2569 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2570 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2571 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2572 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2573 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2574 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2575 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2576 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2577 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2578 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2579 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2580 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2581 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2582 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2583 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2584 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2585 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2586 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2587 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2588 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2589 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2590 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2591 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2592 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2593 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2594 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2595 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2596 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2597 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2598 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2599 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2600 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2601 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2602 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2603 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2604 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2605 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2606 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2607 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2608 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2609 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2610 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2611 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2612 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2613 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2614 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2615 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2616 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2617 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2618 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2619 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2620 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2621 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2622 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2623 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2624 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2625 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2626 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2627 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2628 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2629 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2630 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2631 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2632 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2633 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2634 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2635 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2636 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2637 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2638 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2639 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2640 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2641 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2642 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2643 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2644 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2645 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2646 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2647 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2648 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2649 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2650 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2651 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2652 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2653 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2654 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2655 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2656 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2657 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2658 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2659 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2660 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2661 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2662 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2663 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2664 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2665 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2666 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2667 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2668 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2669 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2670 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2671 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2672 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2673 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2674 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2675 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2676 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2677 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2678 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2679 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2680 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2681 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2682 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2683 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2684 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2685 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2686 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2687 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2688 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2689 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2690 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2691 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2692 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2693 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2694 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2695 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2696 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2697 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2698 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2699 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2700 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2701 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2702 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2703 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2704 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2705 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2706 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2707 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2708 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2709 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2710 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2711 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2712 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2713 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2714 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2715 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2716 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2717 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2718 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2719 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2720 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2721 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2722 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2723 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2724 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2725 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2726 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2727 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2728 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2729 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2730 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2731 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2732 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2733 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2734 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2735 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2736 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2737 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2738 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2739 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2740 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2741 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2742 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2743 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2744 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2745 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2746 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2747 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2748 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2749 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2750 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2751 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2752 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2753 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2754 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2755 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2756 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2757 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2758 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2759 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2760 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2761 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2762 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2763 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2764 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2765 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2766 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2767 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2768 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2769 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2770 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2771 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2772 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2773 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2774 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2775 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2776 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2777 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2778 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2779 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2780 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2781 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2782 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2783 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2784 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2785 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2786 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2787 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2788 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2789 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2790 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2791 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2792 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2793 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2794 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2795 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2796 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2797 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2798 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2799 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2800 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2801 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2802 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2803 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2804 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2805 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2806 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2807 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2808 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2809 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2810 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2811 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2812 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2813 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2814 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2815 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2816 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2817 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2818 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2819 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2820 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2821 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2822 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2823 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2824 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2825 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2826 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2827 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2828 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2829 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2830 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2831 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2832 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2833 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2834 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2835 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2836 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2837 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2838 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2839 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2840 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2841 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2842 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2843 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2844 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2845 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2846 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2847 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2848 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2849 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2850 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2851 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2852 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2853 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2854 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2855 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2856 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2857 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2858 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2859 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2860 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2861 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2862 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2863 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2864 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2865 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2866 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2867 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2868 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2869 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2870 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2871 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2872 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2873 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2874 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2875 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2876 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2877 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2878 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2879 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2880 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2881 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2882 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2883 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2884 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2885 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2886 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2887 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2888 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2889 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2890 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2891 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2892 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2893 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2894 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2895 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2896 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2897 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2898 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2899 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2900 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2901 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2902 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2903 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2904 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2905 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2906 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2907 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2908 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2909 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2910 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2911 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2912 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2913 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2914 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2915 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2916 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2917 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2918 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2919 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2920 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2921 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2922 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2923 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2924 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2925 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2926 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2927 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2928 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2929 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2930 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2931 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2932 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2933 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2934 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2935 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2936 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2937 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2938 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2939 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2940 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2941 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2942 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2943 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2944 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2945 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2946 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2947 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2948 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2949 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2950 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2951 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2952 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2953 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2954 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2955 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2956 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2957 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2958 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2959 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2960 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2961 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2962 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2963 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2964 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2965 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2966 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2967 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2968 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2969 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2970 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2971 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2972 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2973 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2974 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2975 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2976 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2977 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2978 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2979 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2980 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2981 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2982 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2983 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2984 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2985 =>	x"0200017F", -- z: 2 rot: 0 ptr: 383
		2986 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2987 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2988 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2989 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		2990 =>	x"0000027F", -- z: 0 rot: 0 ptr: 639
		others => x"00000000"
	);







begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;